module rock_rom
	(
		input wire clk,
		input wire [5:0] row,
		input wire [5:0] col,
		output reg [11:0] color_data
	);

	(* rom_style = "block" *)

	//signal declaration
	reg [5:0] row_reg;
	reg [5:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @(*) begin







		if(({row_reg, col_reg}>=12'b000000000000) && ({row_reg, col_reg}<12'b000111010101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==12'b000111010101)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=12'b000111010110) && ({row_reg, col_reg}<12'b001000010101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==12'b001000010101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==12'b001000010110)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}==12'b001000010111)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}>=12'b001000011000) && ({row_reg, col_reg}<12'b001000011010)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==12'b001000011010)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}==12'b001000011011)) color_data = 12'b011110101101;

		if(({row_reg, col_reg}>=12'b001000011100) && ({row_reg, col_reg}<12'b001001010100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==12'b001001010100)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}==12'b001001010101)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==12'b001001010110)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==12'b001001010111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==12'b001001011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b001001011001)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==12'b001001011010)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==12'b001001011011)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==12'b001001011100)) color_data = 12'b100010101101;

		if(({row_reg, col_reg}>=12'b001001011101) && ({row_reg, col_reg}<12'b001010010010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==12'b001010010010)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}==12'b001010010011)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==12'b001010010100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=12'b001010010101) && ({row_reg, col_reg}<12'b001010011001)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==12'b001010011001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==12'b001010011010)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==12'b001010011011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==12'b001010011100)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==12'b001010011101)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==12'b001010011110)) color_data = 12'b011010101111;

		if(({row_reg, col_reg}>=12'b001010011111) && ({row_reg, col_reg}<12'b001011010001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==12'b001011010001)) color_data = 12'b011110011100;
		if(({row_reg, col_reg}==12'b001011010010)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}>=12'b001011010011) && ({row_reg, col_reg}<12'b001011010101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==12'b001011010101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b001011010110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=12'b001011010111) && ({row_reg, col_reg}<12'b001011011001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==12'b001011011001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b001011011010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==12'b001011011011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=12'b001011011100) && ({row_reg, col_reg}<12'b001011011110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b001011011110)) color_data = 12'b011110011100;

		if(({row_reg, col_reg}>=12'b001011011111) && ({row_reg, col_reg}<12'b001100010000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==12'b001100010000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==12'b001100010001)) color_data = 12'b100010011010;
		if(({row_reg, col_reg}==12'b001100010010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=12'b001100010011) && ({row_reg, col_reg}<12'b001100010110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==12'b001100010110)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==12'b001100010111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==12'b001100011000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==12'b001100011001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=12'b001100011010) && ({row_reg, col_reg}<12'b001100011101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==12'b001100011101)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==12'b001100011110)) color_data = 12'b011110001000;
		if(({row_reg, col_reg}==12'b001100011111)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=12'b001100100000) && ({row_reg, col_reg}<12'b001101010000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==12'b001101010000)) color_data = 12'b011110011011;
		if(({row_reg, col_reg}==12'b001101010001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=12'b001101010010) && ({row_reg, col_reg}<12'b001101010101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==12'b001101010101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b001101010110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==12'b001101010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b001101011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=12'b001101011001) && ({row_reg, col_reg}<12'b001101011101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==12'b001101011101)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==12'b001101011110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b001101011111)) color_data = 12'b011110011011;
		if(({row_reg, col_reg}==12'b001101100000)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=12'b001101100001) && ({row_reg, col_reg}<12'b001110001111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==12'b001110001111)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==12'b001110010000)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}>=12'b001110010001) && ({row_reg, col_reg}<12'b001110010100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==12'b001110010100)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==12'b001110010101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==12'b001110010110)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==12'b001110010111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=12'b001110011000) && ({row_reg, col_reg}<12'b001110011100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==12'b001110011100)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}>=12'b001110011101) && ({row_reg, col_reg}<12'b001110011111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==12'b001110011111)) color_data = 12'b011110001001;
		if(({row_reg, col_reg}==12'b001110100000)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=12'b001110100001) && ({row_reg, col_reg}<12'b001111001110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==12'b001111001110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==12'b001111001111)) color_data = 12'b011110001010;
		if(({row_reg, col_reg}==12'b001111010000)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==12'b001111010001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b001111010010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=12'b001111010011) && ({row_reg, col_reg}<12'b001111010101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==12'b001111010101)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==12'b001111010110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==12'b001111010111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b001111011000)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=12'b001111011001) && ({row_reg, col_reg}<12'b001111011110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==12'b001111011110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==12'b001111011111)) color_data = 12'b011110001000;
		if(({row_reg, col_reg}==12'b001111100000)) color_data = 12'b011110101101;

		if(({row_reg, col_reg}>=12'b001111100001) && ({row_reg, col_reg}<12'b010000001110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==12'b010000001110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==12'b010000001111)) color_data = 12'b011110011010;
		if(({row_reg, col_reg}==12'b010000010000)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==12'b010000010001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=12'b010000010010) && ({row_reg, col_reg}<12'b010000010100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==12'b010000010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=12'b010000010101) && ({row_reg, col_reg}<12'b010000011110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==12'b010000011110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b010000011111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==12'b010000100000)) color_data = 12'b100010011010;

		if(({row_reg, col_reg}>=12'b010000100001) && ({row_reg, col_reg}<12'b010001001110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==12'b010001001110)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}==12'b010001001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b010001010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=12'b010001010001) && ({row_reg, col_reg}<12'b010001010100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=12'b010001010100) && ({row_reg, col_reg}<12'b010001011100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==12'b010001011100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=12'b010001011101) && ({row_reg, col_reg}<12'b010001011111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==12'b010001011111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==12'b010001100000)) color_data = 12'b100110101011;

		if(({row_reg, col_reg}>=12'b010001100001) && ({row_reg, col_reg}<12'b010010001110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==12'b010010001110)) color_data = 12'b011110011010;
		if(({row_reg, col_reg}==12'b010010001111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=12'b010010010000) && ({row_reg, col_reg}<12'b010010010100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=12'b010010010100) && ({row_reg, col_reg}<12'b010010011010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==12'b010010011010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=12'b010010011011) && ({row_reg, col_reg}<12'b010010011111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==12'b010010011111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==12'b010010100000)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}>=12'b010010100001) && ({row_reg, col_reg}<12'b010010100100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=12'b010010100100) && ({row_reg, col_reg}<12'b010010101000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==12'b010010101000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==12'b010010101001)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=12'b010010101010) && ({row_reg, col_reg}<12'b010011001101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==12'b010011001101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==12'b010011001110)) color_data = 12'b011110001001;
		if(({row_reg, col_reg}>=12'b010011001111) && ({row_reg, col_reg}<12'b010011010100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=12'b010011010100) && ({row_reg, col_reg}<12'b010011011010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=12'b010011011010) && ({row_reg, col_reg}<12'b010011011111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==12'b010011011111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==12'b010011100000)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}>=12'b010011100001) && ({row_reg, col_reg}<12'b010011100011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==12'b010011100011)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==12'b010011100100)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==12'b010011100101)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==12'b010011100110)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==12'b010011100111)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}==12'b010011101000)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=12'b010011101001) && ({row_reg, col_reg}<12'b010100001010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=12'b010100001010) && ({row_reg, col_reg}<12'b010100001100)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==12'b010100001100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==12'b010100001101)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}==12'b010100001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=12'b010100001111) && ({row_reg, col_reg}<12'b010100010100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=12'b010100010100) && ({row_reg, col_reg}<12'b010100011001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=12'b010100011001) && ({row_reg, col_reg}<12'b010100011111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==12'b010100011111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==12'b010100100000)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==12'b010100100001)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==12'b010100100010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==12'b010100100011)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==12'b010100100100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==12'b010100100101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=12'b010100100110) && ({row_reg, col_reg}<12'b010100101000)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==12'b010100101000)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}==12'b010100101001)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=12'b010100101010) && ({row_reg, col_reg}<12'b010101001010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=12'b010101001010) && ({row_reg, col_reg}<12'b010101001100)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==12'b010101001100)) color_data = 12'b011111001110;
		if(({row_reg, col_reg}==12'b010101001101)) color_data = 12'b100111001101;
		if(({row_reg, col_reg}==12'b010101001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=12'b010101001111) && ({row_reg, col_reg}<12'b010101010100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==12'b010101010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b010101010101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b010101010110)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==12'b010101010111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==12'b010101011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=12'b010101011001) && ({row_reg, col_reg}<12'b010101011011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=12'b010101011011) && ({row_reg, col_reg}<12'b010101011101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==12'b010101011101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==12'b010101011110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b010101011111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==12'b010101100000)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==12'b010101100001)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==12'b010101100010)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==12'b010101100011)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==12'b010101100100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b010101100101)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==12'b010101100110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b010101100111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b010101101000)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==12'b010101101001)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}==12'b010101101010)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=12'b010101101011) && ({row_reg, col_reg}<12'b010110001001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=12'b010110001001) && ({row_reg, col_reg}<12'b010110001011)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}==12'b010110001011)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}==12'b010110001100)) color_data = 12'b010010111101;
		if(({row_reg, col_reg}==12'b010110001101)) color_data = 12'b011110111100;
		if(({row_reg, col_reg}==12'b010110001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=12'b010110001111) && ({row_reg, col_reg}<12'b010110010100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==12'b010110010100)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==12'b010110010101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=12'b010110010110) && ({row_reg, col_reg}<12'b010110011000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=12'b010110011000) && ({row_reg, col_reg}<12'b010110011010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==12'b010110011010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b010110011011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==12'b010110011100)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==12'b010110011101)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==12'b010110011110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==12'b010110011111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==12'b010110100000)) color_data = 12'b100010011011;
		if(({row_reg, col_reg}==12'b010110100001)) color_data = 12'b010110001100;
		if(({row_reg, col_reg}==12'b010110100010)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==12'b010110100011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b010110100100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==12'b010110100101)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==12'b010110100110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==12'b010110100111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b010110101000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==12'b010110101001)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==12'b010110101010)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}==12'b010110101011)) color_data = 12'b011110101101;

		if(({row_reg, col_reg}>=12'b010110101100) && ({row_reg, col_reg}<12'b010111000111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==12'b010111000111)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==12'b010111001000)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==12'b010111001001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b010111001010)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==12'b010111001011)) color_data = 12'b100111001100;
		if(({row_reg, col_reg}==12'b010111001100)) color_data = 12'b011011001101;
		if(({row_reg, col_reg}==12'b010111001101)) color_data = 12'b100011001101;
		if(({row_reg, col_reg}==12'b010111001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=12'b010111001111) && ({row_reg, col_reg}<12'b010111010011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==12'b010111010011)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==12'b010111010100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==12'b010111010101)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==12'b010111010110)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==12'b010111010111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==12'b010111011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b010111011001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=12'b010111011010) && ({row_reg, col_reg}<12'b010111011100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==12'b010111011100)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=12'b010111011101) && ({row_reg, col_reg}<12'b010111011111)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==12'b010111011111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b010111100000)) color_data = 12'b011110111101;
		if(({row_reg, col_reg}==12'b010111100001)) color_data = 12'b011010001011;
		if(({row_reg, col_reg}==12'b010111100010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b010111100011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==12'b010111100100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==12'b010111100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b010111100110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==12'b010111100111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==12'b010111101000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=12'b010111101001) && ({row_reg, col_reg}<12'b010111101011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b010111101011)) color_data = 12'b011110001010;
		if(({row_reg, col_reg}==12'b010111101100)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=12'b010111101101) && ({row_reg, col_reg}<12'b011000000100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==12'b011000000100)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=12'b011000000101) && ({row_reg, col_reg}<12'b011000000111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==12'b011000000111)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==12'b011000001000)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==12'b011000001001)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==12'b011000001010)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==12'b011000001011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b011000001100)) color_data = 12'b100110111100;
		if(({row_reg, col_reg}==12'b011000001101)) color_data = 12'b010110011101;
		if(({row_reg, col_reg}==12'b011000001110)) color_data = 12'b011110011011;
		if(({row_reg, col_reg}==12'b011000001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b011000010000)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==12'b011000010001)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==12'b011000010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b011000010011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==12'b011000010100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==12'b011000010101)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==12'b011000010110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b011000010111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b011000011000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=12'b011000011001) && ({row_reg, col_reg}<12'b011000011011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==12'b011000011011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b011000011100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b011000011101)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==12'b011000011110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==12'b011000011111)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==12'b011000100000)) color_data = 12'b011010011011;
		if(({row_reg, col_reg}==12'b011000100001)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==12'b011000100010)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==12'b011000100011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b011000100100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==12'b011000100101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==12'b011000100110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==12'b011000100111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=12'b011000101000) && ({row_reg, col_reg}<12'b011000101010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==12'b011000101010)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==12'b011000101011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b011000101100)) color_data = 12'b011110101101;

		if(({row_reg, col_reg}>=12'b011000101101) && ({row_reg, col_reg}<12'b011001000110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==12'b011001000110)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==12'b011001000111)) color_data = 12'b011110011011;
		if(({row_reg, col_reg}==12'b011001001000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b011001001001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==12'b011001001010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b011001001011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b011001001100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b011001001101)) color_data = 12'b100111001101;
		if(({row_reg, col_reg}==12'b011001001110)) color_data = 12'b010110101101;
		if(({row_reg, col_reg}==12'b011001001111)) color_data = 12'b011010001011;
		if(({row_reg, col_reg}==12'b011001010000)) color_data = 12'b100010011010;
		if(({row_reg, col_reg}==12'b011001010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=12'b011001010010) && ({row_reg, col_reg}<12'b011001010101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==12'b011001010101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=12'b011001010110) && ({row_reg, col_reg}<12'b011001011000)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==12'b011001011000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==12'b011001011001)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==12'b011001011010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b011001011011)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==12'b011001011100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==12'b011001011101)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==12'b011001011110)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==12'b011001011111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b011001100000)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==12'b011001100001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==12'b011001100010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b011001100011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==12'b011001100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b011001100101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==12'b011001100110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b011001100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b011001101000)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==12'b011001101001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b011001101010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==12'b011001101011)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==12'b011001101100)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==12'b011001101101)) color_data = 12'b011110011101;

		if(({row_reg, col_reg}>=12'b011001101110) && ({row_reg, col_reg}<12'b011010000100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=12'b011010000100) && ({row_reg, col_reg}<12'b011010000110)) color_data = 12'b011111001110;
		if(({row_reg, col_reg}==12'b011010000110)) color_data = 12'b011010101100;
		if(({row_reg, col_reg}==12'b011010000111)) color_data = 12'b100110001001;
		if(({row_reg, col_reg}==12'b011010001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b011010001001)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==12'b011010001010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==12'b011010001011)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==12'b011010001100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b011010001101)) color_data = 12'b100110101001;
		if(({row_reg, col_reg}==12'b011010001110)) color_data = 12'b011111001101;
		if(({row_reg, col_reg}==12'b011010001111)) color_data = 12'b001110011101;
		if(({row_reg, col_reg}==12'b011010010000)) color_data = 12'b010110101101;
		if(({row_reg, col_reg}==12'b011010010001)) color_data = 12'b100111001100;
		if(({row_reg, col_reg}==12'b011010010010)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==12'b011010010011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==12'b011010010100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b011010010101)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==12'b011010010110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==12'b011010010111)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==12'b011010011000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==12'b011010011001)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==12'b011010011010)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==12'b011010011011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b011010011100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==12'b011010011101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==12'b011010011110)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==12'b011010011111)) color_data = 12'b100110001001;
		if(({row_reg, col_reg}>=12'b011010100000) && ({row_reg, col_reg}<12'b011010100010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b011010100010)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==12'b011010100011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==12'b011010100100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=12'b011010100101) && ({row_reg, col_reg}<12'b011010100111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==12'b011010100111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b011010101000)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==12'b011010101001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==12'b011010101010)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==12'b011010101011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==12'b011010101100)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==12'b011010101101)) color_data = 12'b011110001001;
		if(({row_reg, col_reg}==12'b011010101110)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=12'b011010101111) && ({row_reg, col_reg}<12'b011011000000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==12'b011011000000)) color_data = 12'b011110111110;
		if(({row_reg, col_reg}>=12'b011011000001) && ({row_reg, col_reg}<12'b011011000011)) color_data = 12'b011111011110;
		if(({row_reg, col_reg}==12'b011011000011)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==12'b011011000100)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==12'b011011000101)) color_data = 12'b011111011110;
		if(({row_reg, col_reg}==12'b011011000110)) color_data = 12'b011010011011;
		if(({row_reg, col_reg}==12'b011011000111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b011011001000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==12'b011011001001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b011011001010)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==12'b011011001011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==12'b011011001100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b011011001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b011011001110)) color_data = 12'b011110101011;
		if(({row_reg, col_reg}==12'b011011001111)) color_data = 12'b010010011110;
		if(({row_reg, col_reg}==12'b011011010000)) color_data = 12'b010110101101;
		if(({row_reg, col_reg}==12'b011011010001)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==12'b011011010010)) color_data = 12'b010101111001;
		if(({row_reg, col_reg}==12'b011011010011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b011011010100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==12'b011011010101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==12'b011011010110)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==12'b011011010111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b011011011000)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==12'b011011011001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b011011011010)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==12'b011011011011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==12'b011011011100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b011011011101)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==12'b011011011110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==12'b011011011111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b011011100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b011011100001)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==12'b011011100010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b011011100011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==12'b011011100100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=12'b011011100101) && ({row_reg, col_reg}<12'b011011101010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==12'b011011101010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b011011101011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b011011101100)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==12'b011011101101)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==12'b011011101110)) color_data = 12'b011110011100;

		if(({row_reg, col_reg}>=12'b011011101111) && ({row_reg, col_reg}<12'b011100000000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==12'b011100000000)) color_data = 12'b011110111110;
		if(({row_reg, col_reg}>=12'b011100000001) && ({row_reg, col_reg}<12'b011100000011)) color_data = 12'b011111001110;
		if(({row_reg, col_reg}==12'b011100000011)) color_data = 12'b010010011101;
		if(({row_reg, col_reg}==12'b011100000100)) color_data = 12'b010010011100;
		if(({row_reg, col_reg}==12'b011100000101)) color_data = 12'b011111011110;
		if(({row_reg, col_reg}==12'b011100000110)) color_data = 12'b010110011010;
		if(({row_reg, col_reg}==12'b011100000111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b011100001000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==12'b011100001001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b011100001010)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==12'b011100001011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==12'b011100001100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==12'b011100001101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==12'b011100001110)) color_data = 12'b010001111010;
		if(({row_reg, col_reg}==12'b011100001111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==12'b011100010000)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}==12'b011100010001)) color_data = 12'b011011001110;
		if(({row_reg, col_reg}==12'b011100010010)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==12'b011100010011)) color_data = 12'b011010001010;
		if(({row_reg, col_reg}==12'b011100010100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b011100010101)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}==12'b011100010110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b011100010111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==12'b011100011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=12'b011100011001) && ({row_reg, col_reg}<12'b011100011011)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==12'b011100011011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==12'b011100011100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=12'b011100011101) && ({row_reg, col_reg}<12'b011100011111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==12'b011100011111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==12'b011100100000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==12'b011100100001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=12'b011100100010) && ({row_reg, col_reg}<12'b011100100100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==12'b011100100100)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==12'b011100100101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=12'b011100100110) && ({row_reg, col_reg}<12'b011100101000)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==12'b011100101000)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==12'b011100101001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==12'b011100101010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=12'b011100101011) && ({row_reg, col_reg}<12'b011100101101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b011100101101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==12'b011100101110)) color_data = 12'b011110001001;
		if(({row_reg, col_reg}==12'b011100101111)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=12'b011100110000) && ({row_reg, col_reg}<12'b011101000000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==12'b011101000000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=12'b011101000001) && ({row_reg, col_reg}<12'b011101000100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==12'b011101000100)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==12'b011101000101)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==12'b011101000110)) color_data = 12'b100011011101;
		if(({row_reg, col_reg}==12'b011101000111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b011101001000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==12'b011101001001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=12'b011101001010) && ({row_reg, col_reg}<12'b011101001110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==12'b011101001110)) color_data = 12'b010001101001;
		if(({row_reg, col_reg}==12'b011101001111)) color_data = 12'b010110111110;
		if(({row_reg, col_reg}==12'b011101010000)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==12'b011101010001)) color_data = 12'b010110111101;
		if(({row_reg, col_reg}==12'b011101010010)) color_data = 12'b100011001110;
		if(({row_reg, col_reg}==12'b011101010011)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==12'b011101010100)) color_data = 12'b100010011011;
		if(({row_reg, col_reg}==12'b011101010101)) color_data = 12'b010001111100;
		if(({row_reg, col_reg}==12'b011101010110)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==12'b011101010111)) color_data = 12'b010101101000;
		if(({row_reg, col_reg}==12'b011101011000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==12'b011101011001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==12'b011101011010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=12'b011101011011) && ({row_reg, col_reg}<12'b011101100000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==12'b011101100000)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==12'b011101100001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=12'b011101100010) && ({row_reg, col_reg}<12'b011101100100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=12'b011101100100) && ({row_reg, col_reg}<12'b011101101000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=12'b011101101000) && ({row_reg, col_reg}<12'b011101101101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==12'b011101101101)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==12'b011101101110)) color_data = 12'b100010101010;
		if(({row_reg, col_reg}==12'b011101101111)) color_data = 12'b100011011111;
		if(({row_reg, col_reg}==12'b011101110000)) color_data = 12'b011010111110;

		if(({row_reg, col_reg}==12'b011101110001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==12'b011110000000)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}>=12'b011110000001) && ({row_reg, col_reg}<12'b011110000100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==12'b011110000100)) color_data = 12'b011111011110;
		if(({row_reg, col_reg}==12'b011110000101)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==12'b011110000110)) color_data = 12'b011111011110;
		if(({row_reg, col_reg}==12'b011110000111)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}==12'b011110001000)) color_data = 12'b010101100111;
		if(({row_reg, col_reg}>=12'b011110001001) && ({row_reg, col_reg}<12'b011110001100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==12'b011110001100)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==12'b011110001101)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==12'b011110001110)) color_data = 12'b010001111011;
		if(({row_reg, col_reg}==12'b011110001111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==12'b011110010000)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==12'b011110010001)) color_data = 12'b100111001110;
		if(({row_reg, col_reg}==12'b011110010010)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==12'b011110010011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==12'b011110010100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==12'b011110010101)) color_data = 12'b011110011100;
		if(({row_reg, col_reg}==12'b011110010110)) color_data = 12'b010010011101;
		if(({row_reg, col_reg}==12'b011110010111)) color_data = 12'b010110101101;
		if(({row_reg, col_reg}==12'b011110011000)) color_data = 12'b010101111000;
		if(({row_reg, col_reg}>=12'b011110011001) && ({row_reg, col_reg}<12'b011110011101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==12'b011110011101)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==12'b011110011110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==12'b011110011111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==12'b011110100000)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}==12'b011110100001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=12'b011110100010) && ({row_reg, col_reg}<12'b011110100101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=12'b011110100101) && ({row_reg, col_reg}<12'b011110101000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==12'b011110101000)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=12'b011110101001) && ({row_reg, col_reg}<12'b011110101101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==12'b011110101101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b011110101110)) color_data = 12'b100011001100;
		if(({row_reg, col_reg}==12'b011110101111)) color_data = 12'b100011011110;
		if(({row_reg, col_reg}==12'b011110110000)) color_data = 12'b011111001110;

		if(({row_reg, col_reg}==12'b011110110001)) color_data = 12'b011110111110;
		if(({row_reg, col_reg}==12'b011111000000)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}==12'b011111000001)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==12'b011111000010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==12'b011111000011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==12'b011111000100)) color_data = 12'b010010011101;
		if(({row_reg, col_reg}==12'b011111000101)) color_data = 12'b011111001110;
		if(({row_reg, col_reg}==12'b011111000110)) color_data = 12'b010010101101;
		if(({row_reg, col_reg}==12'b011111000111)) color_data = 12'b010110101101;
		if(({row_reg, col_reg}==12'b011111001000)) color_data = 12'b011010101100;
		if(({row_reg, col_reg}==12'b011111001001)) color_data = 12'b011010001001;
		if(({row_reg, col_reg}==12'b011111001010)) color_data = 12'b011110011001;
		if(({row_reg, col_reg}==12'b011111001011)) color_data = 12'b011010001001;
		if(({row_reg, col_reg}==12'b011111001100)) color_data = 12'b011110011001;
		if(({row_reg, col_reg}==12'b011111001101)) color_data = 12'b011111001100;
		if(({row_reg, col_reg}==12'b011111001110)) color_data = 12'b011011011110;
		if(({row_reg, col_reg}==12'b011111001111)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==12'b011111010000)) color_data = 12'b010010011101;
		if(({row_reg, col_reg}==12'b011111010001)) color_data = 12'b101010111011;
		if(({row_reg, col_reg}==12'b011111010010)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==12'b011111010011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==12'b011111010100)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==12'b011111010101)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==12'b011111010110)) color_data = 12'b101011011100;
		if(({row_reg, col_reg}==12'b011111010111)) color_data = 12'b011011001110;
		if(({row_reg, col_reg}==12'b011111011000)) color_data = 12'b010110101101;
		if(({row_reg, col_reg}==12'b011111011001)) color_data = 12'b010110001001;
		if(({row_reg, col_reg}==12'b011111011010)) color_data = 12'b011010011001;
		if(({row_reg, col_reg}==12'b011111011011)) color_data = 12'b010101101001;
		if(({row_reg, col_reg}==12'b011111011100)) color_data = 12'b011010011001;
		if(({row_reg, col_reg}==12'b011111011101)) color_data = 12'b100111001011;
		if(({row_reg, col_reg}==12'b011111011110)) color_data = 12'b101011001100;
		if(({row_reg, col_reg}==12'b011111011111)) color_data = 12'b011010011100;
		if(({row_reg, col_reg}==12'b011111100000)) color_data = 12'b001101111011;
		if(({row_reg, col_reg}==12'b011111100001)) color_data = 12'b010101101000;
		if(({row_reg, col_reg}==12'b011111100010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=12'b011111100011) && ({row_reg, col_reg}<12'b011111100110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==12'b011111100110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=12'b011111100111) && ({row_reg, col_reg}<12'b011111101100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==12'b011111101100)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==12'b011111101101)) color_data = 12'b011110101010;
		if(({row_reg, col_reg}==12'b011111101110)) color_data = 12'b011111101111;
		if(({row_reg, col_reg}==12'b011111101111)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==12'b011111110000)) color_data = 12'b011010111110;

		if(({row_reg, col_reg}>=12'b011111110001) && ({row_reg, col_reg}<12'b100000000001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==12'b100000000001)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==12'b100000000010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==12'b100000000011)) color_data = 12'b010010011101;
		if(({row_reg, col_reg}>=12'b100000000100) && ({row_reg, col_reg}<12'b100000000110)) color_data = 12'b010010001110;
		if(({row_reg, col_reg}==12'b100000000110)) color_data = 12'b010010101110;
		if(({row_reg, col_reg}==12'b100000000111)) color_data = 12'b010010101101;
		if(({row_reg, col_reg}==12'b100000001000)) color_data = 12'b010110101101;
		if(({row_reg, col_reg}==12'b100000001001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==12'b100000001010)) color_data = 12'b010110101101;
		if(({row_reg, col_reg}==12'b100000001011)) color_data = 12'b011111101111;
		if(({row_reg, col_reg}==12'b100000001100)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}>=12'b100000001101) && ({row_reg, col_reg}<12'b100000001111)) color_data = 12'b010010101101;
		if(({row_reg, col_reg}>=12'b100000001111) && ({row_reg, col_reg}<12'b100000010001)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}==12'b100000010001)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==12'b100000010010)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==12'b100000010011)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==12'b100000010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==12'b100000010101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==12'b100000010110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==12'b100000010111)) color_data = 12'b011111001101;
		if(({row_reg, col_reg}==12'b100000011000)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==12'b100000011001)) color_data = 12'b011011001110;
		if(({row_reg, col_reg}==12'b100000011010)) color_data = 12'b001110011101;
		if(({row_reg, col_reg}==12'b100000011011)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==12'b100000011100)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}==12'b100000011101)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==12'b100000011110)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==12'b100000011111)) color_data = 12'b011011001110;
		if(({row_reg, col_reg}==12'b100000100000)) color_data = 12'b011011011111;
		if(({row_reg, col_reg}==12'b100000100001)) color_data = 12'b100011011110;
		if(({row_reg, col_reg}==12'b100000100010)) color_data = 12'b011110011000;
		if(({row_reg, col_reg}==12'b100000100011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b100000100100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==12'b100000100101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b100000100110)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}>=12'b100000100111) && ({row_reg, col_reg}<12'b100000101010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==12'b100000101010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==12'b100000101011)) color_data = 12'b010101111001;
		if(({row_reg, col_reg}==12'b100000101100)) color_data = 12'b100011011101;
		if(({row_reg, col_reg}==12'b100000101101)) color_data = 12'b011011001110;
		if(({row_reg, col_reg}==12'b100000101110)) color_data = 12'b010110111101;
		if(({row_reg, col_reg}==12'b100000101111)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==12'b100000110000)) color_data = 12'b010110101101;

		if(({row_reg, col_reg}>=12'b100000110001) && ({row_reg, col_reg}<12'b100001000011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==12'b100001000011)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}>=12'b100001000100) && ({row_reg, col_reg}<12'b100001001000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==12'b100001001000)) color_data = 12'b010010001110;
		if(({row_reg, col_reg}==12'b100001001001)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}==12'b100001001010)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}==12'b100001001011)) color_data = 12'b010010101100;
		if(({row_reg, col_reg}==12'b100001001100)) color_data = 12'b001110011101;
		if(({row_reg, col_reg}>=12'b100001001101) && ({row_reg, col_reg}<12'b100001001111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==12'b100001001111)) color_data = 12'b001110011100;
		if(({row_reg, col_reg}==12'b100001010000)) color_data = 12'b011011001101;
		if(({row_reg, col_reg}==12'b100001010001)) color_data = 12'b011110001001;
		if(({row_reg, col_reg}==12'b100001010010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==12'b100001010011)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=12'b100001010100) && ({row_reg, col_reg}<12'b100001010110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==12'b100001010110)) color_data = 12'b010101111010;
		if(({row_reg, col_reg}==12'b100001010111)) color_data = 12'b010010011101;
		if(({row_reg, col_reg}==12'b100001011000)) color_data = 12'b001110011101;
		if(({row_reg, col_reg}==12'b100001011001)) color_data = 12'b010110101101;
		if(({row_reg, col_reg}==12'b100001011010)) color_data = 12'b010110111110;
		if(({row_reg, col_reg}==12'b100001011011)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==12'b100001011100)) color_data = 12'b011011011110;
		if(({row_reg, col_reg}==12'b100001011101)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==12'b100001011110)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==12'b100001011111)) color_data = 12'b010110111101;
		if(({row_reg, col_reg}==12'b100001100000)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==12'b100001100001)) color_data = 12'b011011011110;
		if(({row_reg, col_reg}==12'b100001100010)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}==12'b100001100011)) color_data = 12'b100111011101;
		if(({row_reg, col_reg}==12'b100001100100)) color_data = 12'b100011001101;
		if(({row_reg, col_reg}>=12'b100001100101) && ({row_reg, col_reg}<12'b100001100111)) color_data = 12'b010001111011;
		if(({row_reg, col_reg}==12'b100001100111)) color_data = 12'b001101111011;
		if(({row_reg, col_reg}==12'b100001101000)) color_data = 12'b011010101100;
		if(({row_reg, col_reg}==12'b100001101001)) color_data = 12'b100111011101;
		if(({row_reg, col_reg}==12'b100001101010)) color_data = 12'b100011011101;
		if(({row_reg, col_reg}==12'b100001101011)) color_data = 12'b011111011110;
		if(({row_reg, col_reg}>=12'b100001101100) && ({row_reg, col_reg}<12'b100001101110)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==12'b100001101110)) color_data = 12'b011111001110;
		if(({row_reg, col_reg}==12'b100001101111)) color_data = 12'b010110101101;
		if(({row_reg, col_reg}==12'b100001110000)) color_data = 12'b010110011101;

		if(({row_reg, col_reg}>=12'b100001110001) && ({row_reg, col_reg}<12'b100010000100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==12'b100010000100)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}>=12'b100010000101) && ({row_reg, col_reg}<12'b100010000111)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==12'b100010000111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==12'b100010001000)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==12'b100010001001)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}==12'b100010001010)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}>=12'b100010001011) && ({row_reg, col_reg}<12'b100010001101)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}==12'b100010001101)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==12'b100010001110)) color_data = 12'b011111101111;
		if(({row_reg, col_reg}==12'b100010001111)) color_data = 12'b011011011110;
		if(({row_reg, col_reg}==12'b100010010000)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}==12'b100010010001)) color_data = 12'b010110011011;
		if(({row_reg, col_reg}==12'b100010010010)) color_data = 12'b011001111000;
		if(({row_reg, col_reg}>=12'b100010010011) && ({row_reg, col_reg}<12'b100010010101)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==12'b100010010101)) color_data = 12'b010001101010;
		if(({row_reg, col_reg}==12'b100010010110)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==12'b100010010111)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==12'b100010011000)) color_data = 12'b001001101101;
		if(({row_reg, col_reg}==12'b100010011001)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==12'b100010011010)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==12'b100010011011)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==12'b100010011100)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==12'b100010011101)) color_data = 12'b011111011110;
		if(({row_reg, col_reg}==12'b100010011110)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==12'b100010011111)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}==12'b100010100000)) color_data = 12'b011011001110;
		if(({row_reg, col_reg}==12'b100010100001)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==12'b100010100010)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==12'b100010100011)) color_data = 12'b001110011101;
		if(({row_reg, col_reg}>=12'b100010100100) && ({row_reg, col_reg}<12'b100010100110)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}>=12'b100010100110) && ({row_reg, col_reg}<12'b100010101000)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==12'b100010101000)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==12'b100010101001)) color_data = 12'b011110111110;
		if(({row_reg, col_reg}==12'b100010101010)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}>=12'b100010101011) && ({row_reg, col_reg}<12'b100010101110)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==12'b100010101110)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}>=12'b100010101111) && ({row_reg, col_reg}<12'b100010110001)) color_data = 12'b011010101110;

		if(({row_reg, col_reg}==12'b100010110001)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=12'b100011000000) && ({row_reg, col_reg}<12'b100011000101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==12'b100011000101)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==12'b100011000110)) color_data = 12'b010010011110;
		if(({row_reg, col_reg}==12'b100011000111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==12'b100011001000)) color_data = 12'b010010001110;
		if(({row_reg, col_reg}>=12'b100011001001) && ({row_reg, col_reg}<12'b100011001100)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==12'b100011001100)) color_data = 12'b010010011101;
		if(({row_reg, col_reg}==12'b100011001101)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==12'b100011001110)) color_data = 12'b011011001110;
		if(({row_reg, col_reg}==12'b100011001111)) color_data = 12'b010010101101;
		if(({row_reg, col_reg}==12'b100011010000)) color_data = 12'b010110101101;
		if(({row_reg, col_reg}==12'b100011010001)) color_data = 12'b011111011110;
		if(({row_reg, col_reg}==12'b100011010010)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}>=12'b100011010011) && ({row_reg, col_reg}<12'b100011010101)) color_data = 12'b011011001101;
		if(({row_reg, col_reg}==12'b100011010101)) color_data = 12'b010010011101;
		if(({row_reg, col_reg}==12'b100011010110)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==12'b100011010111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==12'b100011011000)) color_data = 12'b010010101101;
		if(({row_reg, col_reg}==12'b100011011001)) color_data = 12'b010010011101;
		if(({row_reg, col_reg}>=12'b100011011010) && ({row_reg, col_reg}<12'b100011011100)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==12'b100011011100)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==12'b100011011101)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}==12'b100011011110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==12'b100011011111)) color_data = 12'b010010011101;
		if(({row_reg, col_reg}>=12'b100011100000) && ({row_reg, col_reg}<12'b100011100010)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}==12'b100011100010)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==12'b100011100011)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==12'b100011100100)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}>=12'b100011100101) && ({row_reg, col_reg}<12'b100011101011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==12'b100011101011)) color_data = 12'b010010001110;
		if(({row_reg, col_reg}==12'b100011101100)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==12'b100011101101)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}==12'b100011101110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=12'b100011101111) && ({row_reg, col_reg}<12'b100011110001)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=12'b100011110001) && ({row_reg, col_reg}<12'b100100000100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==12'b100100000100)) color_data = 12'b010010011110;
		if(({row_reg, col_reg}==12'b100100000101)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==12'b100100000110)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==12'b100100000111)) color_data = 12'b010010001110;
		if(({row_reg, col_reg}==12'b100100001000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=12'b100100001001) && ({row_reg, col_reg}<12'b100100001011)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==12'b100100001011)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==12'b100100001100)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==12'b100100001101)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}==12'b100100001110)) color_data = 12'b010110101101;
		if(({row_reg, col_reg}==12'b100100001111)) color_data = 12'b010110111110;
		if(({row_reg, col_reg}==12'b100100010000)) color_data = 12'b010110111101;
		if(({row_reg, col_reg}==12'b100100010001)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==12'b100100010010)) color_data = 12'b010110111101;
		if(({row_reg, col_reg}==12'b100100010011)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==12'b100100010100)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==12'b100100010101)) color_data = 12'b011111011110;
		if(({row_reg, col_reg}==12'b100100010110)) color_data = 12'b010110111101;
		if(({row_reg, col_reg}==12'b100100010111)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==12'b100100011000)) color_data = 12'b010110111101;
		if(({row_reg, col_reg}==12'b100100011001)) color_data = 12'b011111001110;
		if(({row_reg, col_reg}>=12'b100100011010) && ({row_reg, col_reg}<12'b100100011100)) color_data = 12'b010110011110;

		if(({row_reg, col_reg}>=12'b100100011100) && ({row_reg, col_reg}<12'b100101000100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==12'b100101000100)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}>=12'b100101000101) && ({row_reg, col_reg}<12'b100101000111)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==12'b100101000111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==12'b100101001000)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==12'b100101001001)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}>=12'b100101001010) && ({row_reg, col_reg}<12'b100101010001)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==12'b100101010001)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==12'b100101010010)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==12'b100101010011)) color_data = 12'b010010101101;
		if(({row_reg, col_reg}==12'b100101010100)) color_data = 12'b010110101101;
		if(({row_reg, col_reg}==12'b100101010101)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==12'b100101010110)) color_data = 12'b010010011101;
		if(({row_reg, col_reg}==12'b100101010111)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==12'b100101011000)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}==12'b100101011001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=12'b100101011010) && ({row_reg, col_reg}<12'b100101011100)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=12'b100101011100) && ({row_reg, col_reg}<12'b100110000110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==12'b100110000110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==12'b100110000111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==12'b100110001000)) color_data = 12'b011110111110;
		if(({row_reg, col_reg}==12'b100110001001)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}==12'b100110001010)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==12'b100110001011)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==12'b100110001100)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==12'b100110001101)) color_data = 12'b010110101110;
		if(({row_reg, col_reg}==12'b100110001110)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}==12'b100110001111)) color_data = 12'b010010011101;
		if(({row_reg, col_reg}==12'b100110010000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==12'b100110010001)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==12'b100110010010)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==12'b100110010011)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==12'b100110010100)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}>=12'b100110010101) && ({row_reg, col_reg}<12'b100110011000)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==12'b100110011000)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=12'b100110011001) && ({row_reg, col_reg}<12'b100111001101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==12'b100111001101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=12'b100111001110) && ({row_reg, col_reg}<12'b100111010000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==12'b100111010000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=12'b100111010001) && ({row_reg, col_reg}<12'b100111010101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=12'b100111010101) && ({row_reg, col_reg}<12'b100111011000)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=12'b100111011000) && ({row_reg, col_reg}<12'b101000001100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==12'b101000001100)) color_data = 12'b011110101110;










		if(({row_reg, col_reg}>=12'b101000001101) && ({row_reg, col_reg}<=12'b110001110001)) color_data = 12'b011010101110;
	end
endmodule