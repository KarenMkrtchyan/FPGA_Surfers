module rock_rom
	(
		input wire clk,
		input wire [8:0] row,
		input wire [8:0] col,
		output reg [11:0] color_data
	);

	(* rom_style = "block" *)

	//signal declaration
	reg [8:0] row_reg;
	reg [8:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @(*) begin
































		if(({row_reg, col_reg}>=18'b000000000000000000) && ({row_reg, col_reg}<18'b000100000010011111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b000100000010011111)) color_data = 12'b011110101110;



		if(({row_reg, col_reg}>=18'b000100000010100000) && ({row_reg, col_reg}<18'b000100011001110100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b000100011001110100) && ({row_reg, col_reg}<18'b000100011001110110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b000100011001110110) && ({row_reg, col_reg}<18'b000100011010000111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b000100011010000111) && ({row_reg, col_reg}<18'b000100011010001001)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b000100011010001001) && ({row_reg, col_reg}<18'b000100011010001111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b000100011010001111)) color_data = 12'b011010101111;

		if(({row_reg, col_reg}>=18'b000100011010010000) && ({row_reg, col_reg}<18'b000100100001110001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b000100100001110001) && ({row_reg, col_reg}<18'b000100100001111001)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b000100100001111001) && ({row_reg, col_reg}<18'b000100101001110100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b000100101001110100) && ({row_reg, col_reg}<18'b000100101001111010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b000100101001111010)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}>=18'b000100101001111011) && ({row_reg, col_reg}<18'b000100101010000000)) color_data = 12'b011010101111;

		if(({row_reg, col_reg}>=18'b000100101010000000) && ({row_reg, col_reg}<18'b000100110001110110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b000100110001110110) && ({row_reg, col_reg}<18'b000100110001111100)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b000100110001111100) && ({row_reg, col_reg}<18'b000100110010000000)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b000100110010000000) && ({row_reg, col_reg}<18'b000100110010000011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b000100110010000011) && ({row_reg, col_reg}<18'b000100110010001010)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b000100110010001010) && ({row_reg, col_reg}<18'b000100110010010101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b000100110010010101) && ({row_reg, col_reg}<18'b000100110010011000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b000100110010011000) && ({row_reg, col_reg}<18'b000100110010011111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b000100110010011111)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b000100110010100000) && ({row_reg, col_reg}<18'b000100111001110111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b000100111001110111) && ({row_reg, col_reg}<18'b000100111001111101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b000100111001111101) && ({row_reg, col_reg}<18'b000100111010010101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b000100111010010101) && ({row_reg, col_reg}<18'b000100111010011001)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b000100111010011001) && ({row_reg, col_reg}<18'b000100111010011100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b000100111010011100) && ({row_reg, col_reg}<18'b000100111010100000)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b000100111010100000) && ({row_reg, col_reg}<18'b000101000001110111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b000101000001110111) && ({row_reg, col_reg}<18'b000101000001111011)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b000101000001111011) && ({row_reg, col_reg}<18'b000101000001111101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b000101000001111101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b000101000001111110) && ({row_reg, col_reg}<18'b000101000010000010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b000101000010000010) && ({row_reg, col_reg}<18'b000101000010000101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b000101000010000101) && ({row_reg, col_reg}<18'b000101000010011101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b000101000010011101) && ({row_reg, col_reg}<18'b000101000010100000)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b000101000010100000) && ({row_reg, col_reg}<18'b000101001001111010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b000101001001111010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b000101001001111011) && ({row_reg, col_reg}<18'b000101001010010000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b000101001010010000) && ({row_reg, col_reg}<18'b000101001010010011)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b000101001010010011) && ({row_reg, col_reg}<18'b000101001010011111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b000101001010011111)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b000101001010100000) && ({row_reg, col_reg}<18'b000101010001110000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b000101010001110000) && ({row_reg, col_reg}<18'b000101010001111000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b000101010001111000) && ({row_reg, col_reg}<18'b000101010001111010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b000101010001111010) && ({row_reg, col_reg}<18'b000101010001111100)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b000101010001111100) && ({row_reg, col_reg}<18'b000101010010000000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b000101010010000000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b000101010010000001) && ({row_reg, col_reg}<18'b000101010010010000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b000101010010010000) && ({row_reg, col_reg}<18'b000101010010010100)) color_data = 12'b011110101111;

		if(({row_reg, col_reg}>=18'b000101010010010100) && ({row_reg, col_reg}<18'b000101011001110000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b000101011001110000) && ({row_reg, col_reg}<18'b000101011010000110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b000101011010000110) && ({row_reg, col_reg}<18'b000101011010001101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b000101011010001101) && ({row_reg, col_reg}<18'b000101011010010000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b000101011010010000)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}>=18'b000101011010010001) && ({row_reg, col_reg}<18'b000101011010010110)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b000101011010010110) && ({row_reg, col_reg}<18'b000101100001110000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b000101100001110000) && ({row_reg, col_reg}<18'b000101100010001110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b000101100010001110) && ({row_reg, col_reg}<18'b000101100010010000)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b000101100010010000) && ({row_reg, col_reg}<18'b000101100010010111)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b000101100010010111) && ({row_reg, col_reg}<18'b000101101001110000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b000101101001110000) && ({row_reg, col_reg}<18'b000101101001111011)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b000101101001111011) && ({row_reg, col_reg}<18'b000101101010010000)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b000101101010010000)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}>=18'b000101101010010001) && ({row_reg, col_reg}<18'b000101101010010100)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}>=18'b000101101010010100) && ({row_reg, col_reg}<18'b000101101010010111)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b000101101010010111)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b000101101010011000) && ({row_reg, col_reg}<18'b000101110001101111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b000101110001101111)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b000101110001110000) && ({row_reg, col_reg}<18'b000101110001110100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b000101110001110100) && ({row_reg, col_reg}<18'b000101110001111000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b000101110001111000) && ({row_reg, col_reg}<18'b000101110001111011)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b000101110001111011) && ({row_reg, col_reg}<18'b000101110001111101)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}>=18'b000101110001111101) && ({row_reg, col_reg}<18'b000101110010010000)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b000101110010010000)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}>=18'b000101110010010001) && ({row_reg, col_reg}<18'b000101110010010101)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}>=18'b000101110010010101) && ({row_reg, col_reg}<18'b000101110010011000)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b000101110010011000)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b000101110010011001) && ({row_reg, col_reg}<18'b000101111001101110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b000101111001101110) && ({row_reg, col_reg}<18'b000101111001110000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b000101111001110000) && ({row_reg, col_reg}<18'b000101111001110101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b000101111001110101) && ({row_reg, col_reg}<18'b000101111001110111)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b000101111001110111) && ({row_reg, col_reg}<18'b000101111001111010)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b000101111001111010)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}==18'b000101111001111011)) color_data = 12'b100010111101;
		if(({row_reg, col_reg}>=18'b000101111001111100) && ({row_reg, col_reg}<18'b000101111010000011)) color_data = 12'b100110111100;
		if(({row_reg, col_reg}>=18'b000101111010000011) && ({row_reg, col_reg}<18'b000101111010000101)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}>=18'b000101111010000101) && ({row_reg, col_reg}<18'b000101111010010000)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}>=18'b000101111010010000) && ({row_reg, col_reg}<18'b000101111010010010)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}>=18'b000101111010010010) && ({row_reg, col_reg}<18'b000101111010010100)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}>=18'b000101111010010100) && ({row_reg, col_reg}<18'b000101111010010110)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}>=18'b000101111010010110) && ({row_reg, col_reg}<18'b000101111010011000)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b000101111010011000)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b000101111010011001) && ({row_reg, col_reg}<18'b000110000001110100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b000110000001110100) && ({row_reg, col_reg}<18'b000110000001110111)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b000110000001110111) && ({row_reg, col_reg}<18'b000110000001111010)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b000110000001111010)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b000110000001111011)) color_data = 12'b100110111100;
		if(({row_reg, col_reg}==18'b000110000001111100)) color_data = 12'b101010111011;
		if(({row_reg, col_reg}==18'b000110000001111101)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}>=18'b000110000001111110) && ({row_reg, col_reg}<18'b000110000010000000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b000110000010000000) && ({row_reg, col_reg}<18'b000110000010000101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b000110000010000101)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==18'b000110000010000110)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}>=18'b000110000010000111) && ({row_reg, col_reg}<18'b000110000010001010)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==18'b000110000010001010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b000110000010001011)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==18'b000110000010001100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b000110000010001101)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}>=18'b000110000010001110) && ({row_reg, col_reg}<18'b000110000010010000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b000110000010010000) && ({row_reg, col_reg}<18'b000110000010010010)) color_data = 12'b101010101000;
		if(({row_reg, col_reg}==18'b000110000010010010)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b000110000010010011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b000110000010010100)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==18'b000110000010010101)) color_data = 12'b100110011011;
		if(({row_reg, col_reg}==18'b000110000010010110)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b000110000010010111)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}==18'b000110000010011000)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b000110000010011001) && ({row_reg, col_reg}<18'b000110000010011011)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b000110000010011011) && ({row_reg, col_reg}<18'b000110001001110001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b000110001001110001) && ({row_reg, col_reg}<18'b000110001001110101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b000110001001110101) && ({row_reg, col_reg}<18'b000110001001111001)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b000110001001111001) && ({row_reg, col_reg}<18'b000110001001111011)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b000110001001111011)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==18'b000110001001111100)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}>=18'b000110001001111101) && ({row_reg, col_reg}<18'b000110001001111111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b000110001001111111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b000110001010000000) && ({row_reg, col_reg}<18'b000110001010000101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b000110001010000101)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==18'b000110001010000110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b000110001010000111)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}>=18'b000110001010001000) && ({row_reg, col_reg}<18'b000110001010001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b000110001010001111)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}>=18'b000110001010010000) && ({row_reg, col_reg}<18'b000110001010010011)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b000110001010010011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b000110001010010100) && ({row_reg, col_reg}<18'b000110001010010110)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}==18'b000110001010010110)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b000110001010010111)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b000110001010011000)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}==18'b000110001010011001)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b000110001010011010) && ({row_reg, col_reg}<18'b000110001010011100)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b000110001010011100) && ({row_reg, col_reg}<18'b000110010001110000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b000110010001110000) && ({row_reg, col_reg}<18'b000110010001110101)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b000110010001110101) && ({row_reg, col_reg}<18'b000110010001110111)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}>=18'b000110010001110111) && ({row_reg, col_reg}<18'b000110010001111010)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b000110010001111010)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}>=18'b000110010001111011) && ({row_reg, col_reg}<18'b000110010001111101)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b000110010001111101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b000110010001111110) && ({row_reg, col_reg}<18'b000110010010000100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b000110010010000100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b000110010010000101) && ({row_reg, col_reg}<18'b000110010010001010)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}>=18'b000110010010001010) && ({row_reg, col_reg}<18'b000110010010001110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b000110010010001110)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}>=18'b000110010010001111) && ({row_reg, col_reg}<18'b000110010010010100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b000110010010010100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b000110010010010101)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}>=18'b000110010010010110) && ({row_reg, col_reg}<18'b000110010010011000)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}>=18'b000110010010011000) && ({row_reg, col_reg}<18'b000110010010011010)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}>=18'b000110010010011010) && ({row_reg, col_reg}<18'b000110010010011101)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b000110010010011101) && ({row_reg, col_reg}<18'b000110010010011111)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b000110010010011111) && ({row_reg, col_reg}<18'b000110010010101001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b000110010010101001) && ({row_reg, col_reg}<18'b000110010010101011)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b000110010010101011) && ({row_reg, col_reg}<18'b000110011001101101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b000110011001101101) && ({row_reg, col_reg}<18'b000110011001110000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b000110011001110000) && ({row_reg, col_reg}<18'b000110011001110010)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}==18'b000110011001110010)) color_data = 12'b100010111101;
		if(({row_reg, col_reg}>=18'b000110011001110011) && ({row_reg, col_reg}<18'b000110011001110101)) color_data = 12'b100110101101;
		if(({row_reg, col_reg}>=18'b000110011001110101) && ({row_reg, col_reg}<18'b000110011001111001)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==18'b000110011001111001)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}>=18'b000110011001111010) && ({row_reg, col_reg}<18'b000110011001111101)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}>=18'b000110011001111101) && ({row_reg, col_reg}<18'b000110011010010010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b000110011010010010)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b000110011010010011) && ({row_reg, col_reg}<18'b000110011010010101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b000110011010010101)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b000110011010010110)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}==18'b000110011010010111)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==18'b000110011010011000)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b000110011010011001)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}>=18'b000110011010011010) && ({row_reg, col_reg}<18'b000110011010011100)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b000110011010011100)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b000110011010011101) && ({row_reg, col_reg}<18'b000110011010100000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b000110011010100000) && ({row_reg, col_reg}<18'b000110011010101001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b000110011010101001) && ({row_reg, col_reg}<18'b000110011010101011)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b000110011010101011) && ({row_reg, col_reg}<18'b000110100001100000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b000110100001100000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b000110100001100001) && ({row_reg, col_reg}<18'b000110100001101100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b000110100001101100) && ({row_reg, col_reg}<18'b000110100001110000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b000110100001110000)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}>=18'b000110100001110001) && ({row_reg, col_reg}<18'b000110100001110011)) color_data = 12'b100110111101;
		if(({row_reg, col_reg}>=18'b000110100001110011) && ({row_reg, col_reg}<18'b000110100001110110)) color_data = 12'b101010101100;
		if(({row_reg, col_reg}>=18'b000110100001110110) && ({row_reg, col_reg}<18'b000110100001111011)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b000110100001111011)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}>=18'b000110100001111100) && ({row_reg, col_reg}<18'b000110100010010010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b000110100010010010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b000110100010010011) && ({row_reg, col_reg}<18'b000110100010010110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b000110100010010110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b000110100010010111)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b000110100010011000) && ({row_reg, col_reg}<18'b000110100010011010)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==18'b000110100010011010)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}>=18'b000110100010011011) && ({row_reg, col_reg}<18'b000110100010011101)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b000110100010011101)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b000110100010011110) && ({row_reg, col_reg}<18'b000110100010100000)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b000110100010100000) && ({row_reg, col_reg}<18'b000110101001100111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b000110101001100111) && ({row_reg, col_reg}<18'b000110101001101010)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}>=18'b000110101001101010) && ({row_reg, col_reg}<18'b000110101001110000)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b000110101001110000)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}==18'b000110101001110001)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==18'b000110101001110010)) color_data = 12'b101010101100;
		if(({row_reg, col_reg}>=18'b000110101001110011) && ({row_reg, col_reg}<18'b000110101001110111)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}>=18'b000110101001110111) && ({row_reg, col_reg}<18'b000110101001111010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b000110101001111010) && ({row_reg, col_reg}<18'b000110101010010010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b000110101010010010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b000110101010010011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b000110101010010100) && ({row_reg, col_reg}<18'b000110101010010110)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b000110101010010110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b000110101010010111) && ({row_reg, col_reg}<18'b000110101010011001)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b000110101010011001) && ({row_reg, col_reg}<18'b000110101010011011)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==18'b000110101010011011)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b000110101010011100)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b000110101010011101)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}==18'b000110101010011110)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b000110101010011111) && ({row_reg, col_reg}<18'b000110101010100011)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b000110101010100011) && ({row_reg, col_reg}<18'b000110110001100110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b000110110001100110)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}>=18'b000110110001100111) && ({row_reg, col_reg}<18'b000110110001101100)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b000110110001101100)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}>=18'b000110110001101101) && ({row_reg, col_reg}<18'b000110110001110000)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}>=18'b000110110001110000) && ({row_reg, col_reg}<18'b000110110001110010)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}>=18'b000110110001110010) && ({row_reg, col_reg}<18'b000110110001110100)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}>=18'b000110110001110100) && ({row_reg, col_reg}<18'b000110110010010010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b000110110010010010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b000110110010010011)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b000110110010010100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b000110110010010101)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b000110110010010110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b000110110010010111) && ({row_reg, col_reg}<18'b000110110010011001)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b000110110010011001) && ({row_reg, col_reg}<18'b000110110010011011)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==18'b000110110010011011)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b000110110010011100)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}==18'b000110110010011101)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b000110110010011110)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}==18'b000110110010011111)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b000110110010100000) && ({row_reg, col_reg}<18'b000110110010100100)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b000110110010100100) && ({row_reg, col_reg}<18'b000110111001100000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b000110111001100000) && ({row_reg, col_reg}<18'b000110111001100010)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b000110111001100010) && ({row_reg, col_reg}<18'b000110111001100101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b000110111001100101) && ({row_reg, col_reg}<18'b000110111001100111)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b000110111001100111) && ({row_reg, col_reg}<18'b000110111001101010)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}>=18'b000110111001101010) && ({row_reg, col_reg}<18'b000110111001101110)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}>=18'b000110111001101110) && ({row_reg, col_reg}<18'b000110111001110000)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b000110111001110000)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}>=18'b000110111001110001) && ({row_reg, col_reg}<18'b000110111001110011)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}>=18'b000110111001110011) && ({row_reg, col_reg}<18'b000110111010000000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b000110111010000000) && ({row_reg, col_reg}<18'b000110111010000010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b000110111010000010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b000110111010000011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b000110111010000100) && ({row_reg, col_reg}<18'b000110111010001110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b000110111010001110) && ({row_reg, col_reg}<18'b000110111010010010)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b000110111010010010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b000110111010010011) && ({row_reg, col_reg}<18'b000110111010010101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b000110111010010101)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b000110111010010110) && ({row_reg, col_reg}<18'b000110111010011000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b000110111010011000)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b000110111010011001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b000110111010011010) && ({row_reg, col_reg}<18'b000110111010011100)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==18'b000110111010011100)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}>=18'b000110111010011101) && ({row_reg, col_reg}<18'b000110111010100000)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}>=18'b000110111010100000) && ({row_reg, col_reg}<18'b000110111010100011)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b000110111010100011)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b000110111010100100) && ({row_reg, col_reg}<18'b000110111010100110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b000110111010100110) && ({row_reg, col_reg}<18'b000110111010101011)) color_data = 12'b011010101111;

		if(({row_reg, col_reg}>=18'b000110111010101011) && ({row_reg, col_reg}<18'b000111000001100000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b000111000001100000)) color_data = 12'b010110101110;
		if(({row_reg, col_reg}>=18'b000111000001100001) && ({row_reg, col_reg}<18'b000111000001100011)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b000111000001100011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b000111000001100100)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b000111000001100101) && ({row_reg, col_reg}<18'b000111000001100111)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b000111000001100111)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}>=18'b000111000001101000) && ({row_reg, col_reg}<18'b000111000001101011)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}>=18'b000111000001101011) && ({row_reg, col_reg}<18'b000111000001101101)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}>=18'b000111000001101101) && ({row_reg, col_reg}<18'b000111000001110000)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}>=18'b000111000001110000) && ({row_reg, col_reg}<18'b000111000001110010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b000111000001110010) && ({row_reg, col_reg}<18'b000111000010001101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b000111000010001101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b000111000010001110) && ({row_reg, col_reg}<18'b000111000010010010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b000111000010010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b000111000010010011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b000111000010010100) && ({row_reg, col_reg}<18'b000111000010010110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b000111000010010110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b000111000010010111)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==18'b000111000010011000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b000111000010011001) && ({row_reg, col_reg}<18'b000111000010011011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b000111000010011011)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}==18'b000111000010011100)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==18'b000111000010011101)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b000111000010011110)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}==18'b000111000010011111)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b000111000010100000)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b000111000010100001)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}>=18'b000111000010100010) && ({row_reg, col_reg}<18'b000111000010100100)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b000111000010100100)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b000111000010100101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b000111000010100110) && ({row_reg, col_reg}<18'b000111000010101100)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b000111000010101100) && ({row_reg, col_reg}<18'b000111000010101111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b000111000010101111)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b000111000010110000) && ({row_reg, col_reg}<18'b000111001001011110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b000111001001011110) && ({row_reg, col_reg}<18'b000111001001100000)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b000111001001100000)) color_data = 12'b011010111111;
		if(({row_reg, col_reg}==18'b000111001001100001)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b000111001001100010) && ({row_reg, col_reg}<18'b000111001001100100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b000111001001100100)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b000111001001100101)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b000111001001100110)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}>=18'b000111001001100111) && ({row_reg, col_reg}<18'b000111001001101001)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}==18'b000111001001101001)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}>=18'b000111001001101010) && ({row_reg, col_reg}<18'b000111001001101100)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==18'b000111001001101100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b000111001001101101) && ({row_reg, col_reg}<18'b000111001001101111)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}>=18'b000111001001101111) && ({row_reg, col_reg}<18'b000111001001110001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b000111001001110001) && ({row_reg, col_reg}<18'b000111001001111111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b000111001001111111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b000111001010000000) && ({row_reg, col_reg}<18'b000111001010001100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b000111001010001100)) color_data = 12'b110010111011;
		if(({row_reg, col_reg}==18'b000111001010001101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b000111001010001110) && ({row_reg, col_reg}<18'b000111001010010010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b000111001010010010)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b000111001010010011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b000111001010010100) && ({row_reg, col_reg}<18'b000111001010011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b000111001010011000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b000111001010011001)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b000111001010011010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b000111001010011011)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}>=18'b000111001010011100) && ({row_reg, col_reg}<18'b000111001010011110)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}>=18'b000111001010011110) && ({row_reg, col_reg}<18'b000111001010100000)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}>=18'b000111001010100000) && ({row_reg, col_reg}<18'b000111001010100010)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b000111001010100010)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}==18'b000111001010100011)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b000111001010100100)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b000111001010100101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b000111001010100110) && ({row_reg, col_reg}<18'b000111001010101100)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b000111001010101100) && ({row_reg, col_reg}<18'b000111001010101110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b000111001010101110) && ({row_reg, col_reg}<18'b000111001010110000)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b000111001010110000) && ({row_reg, col_reg}<18'b000111010001011100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b000111010001011100)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b000111010001011101) && ({row_reg, col_reg}<18'b000111010001100000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b000111010001100000)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b000111010001100001) && ({row_reg, col_reg}<18'b000111010001100011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b000111010001100011)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b000111010001100100)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b000111010001100101)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}==18'b000111010001100110)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b000111010001100111)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}==18'b000111010001101000)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b000111010001101001)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==18'b000111010001101010)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}==18'b000111010001101011)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==18'b000111010001101100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b000111010001101101) && ({row_reg, col_reg}<18'b000111010010001101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b000111010010001101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b000111010010001110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b000111010010001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b000111010010010000) && ({row_reg, col_reg}<18'b000111010010010010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b000111010010010010)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b000111010010010011)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b000111010010010100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b000111010010010101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b000111010010010110) && ({row_reg, col_reg}<18'b000111010010011100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b000111010010011100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b000111010010011101)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==18'b000111010010011110)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}==18'b000111010010011111)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}>=18'b000111010010100000) && ({row_reg, col_reg}<18'b000111010010100011)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b000111010010100011)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}==18'b000111010010100100)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b000111010010100101) && ({row_reg, col_reg}<18'b000111010010100111)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b000111010010100111) && ({row_reg, col_reg}<18'b000111010010101101)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b000111010010101101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b000111010010101110) && ({row_reg, col_reg}<18'b000111010010110000)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b000111010010110000) && ({row_reg, col_reg}<18'b000111011001100010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b000111011001100010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b000111011001100011) && ({row_reg, col_reg}<18'b000111011001100101)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b000111011001100101)) color_data = 12'b100010011100;
		if(({row_reg, col_reg}==18'b000111011001100110)) color_data = 12'b100010011011;
		if(({row_reg, col_reg}==18'b000111011001100111)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b000111011001101000)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}==18'b000111011001101001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b000111011001101010)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}>=18'b000111011001101011) && ({row_reg, col_reg}<18'b000111011001101101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b000111011001101101) && ({row_reg, col_reg}<18'b000111011001111000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b000111011001111000)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}>=18'b000111011001111001) && ({row_reg, col_reg}<18'b000111011010000100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b000111011010000100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b000111011010000101) && ({row_reg, col_reg}<18'b000111011010001101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b000111011010001101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b000111011010001110)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}>=18'b000111011010001111) && ({row_reg, col_reg}<18'b000111011010010010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b000111011010010010)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b000111011010010011) && ({row_reg, col_reg}<18'b000111011010010111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b000111011010010111) && ({row_reg, col_reg}<18'b000111011010011001)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b000111011010011001) && ({row_reg, col_reg}<18'b000111011010011100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b000111011010011100) && ({row_reg, col_reg}<18'b000111011010011110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b000111011010011110)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==18'b000111011010011111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b000111011010100000)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b000111011010100001)) color_data = 12'b100010011011;
		if(({row_reg, col_reg}>=18'b000111011010100010) && ({row_reg, col_reg}<18'b000111011010100100)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b000111011010100100)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}==18'b000111011010100101)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b000111011010100110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b000111011010100111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b000111011010101000) && ({row_reg, col_reg}<18'b000111011010101011)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b000111011010101011) && ({row_reg, col_reg}<18'b000111011010101110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b000111011010101110)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b000111011010101111) && ({row_reg, col_reg}<18'b000111100001100000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b000111100001100000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b000111100001100001) && ({row_reg, col_reg}<18'b000111100001100011)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b000111100001100011) && ({row_reg, col_reg}<18'b000111100001100101)) color_data = 12'b011010001011;
		if(({row_reg, col_reg}==18'b000111100001100101)) color_data = 12'b011110001010;
		if(({row_reg, col_reg}==18'b000111100001100110)) color_data = 12'b100010001010;
		if(({row_reg, col_reg}==18'b000111100001100111)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}>=18'b000111100001101000) && ({row_reg, col_reg}<18'b000111100001101101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b000111100001101101) && ({row_reg, col_reg}<18'b000111100001110110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b000111100001110110) && ({row_reg, col_reg}<18'b000111100001111000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b000111100001111000) && ({row_reg, col_reg}<18'b000111100010000100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b000111100010000100) && ({row_reg, col_reg}<18'b000111100010000111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b000111100010000111)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b000111100010001000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b000111100010001001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b000111100010001010) && ({row_reg, col_reg}<18'b000111100010001101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b000111100010001101)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b000111100010001110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b000111100010001111) && ({row_reg, col_reg}<18'b000111100010010010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b000111100010010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b000111100010010011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b000111100010010100) && ({row_reg, col_reg}<18'b000111100010010110)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b000111100010010110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b000111100010010111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b000111100010011000) && ({row_reg, col_reg}<18'b000111100010011010)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b000111100010011010)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b000111100010011011)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b000111100010011100) && ({row_reg, col_reg}<18'b000111100010011111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b000111100010011111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b000111100010100000)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b000111100010100001)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}==18'b000111100010100010)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}>=18'b000111100010100011) && ({row_reg, col_reg}<18'b000111100010100101)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b000111100010100101)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}==18'b000111100010100110)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b000111100010100111) && ({row_reg, col_reg}<18'b000111100010101010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b000111100010101010) && ({row_reg, col_reg}<18'b000111100010101110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b000111100010101110)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b000111100010101111) && ({row_reg, col_reg}<18'b000111101001011110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b000111101001011110) && ({row_reg, col_reg}<18'b000111101001100000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b000111101001100000) && ({row_reg, col_reg}<18'b000111101001100010)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b000111101001100010)) color_data = 12'b011110011100;
		if(({row_reg, col_reg}>=18'b000111101001100011) && ({row_reg, col_reg}<18'b000111101001100101)) color_data = 12'b011010001010;
		if(({row_reg, col_reg}==18'b000111101001100101)) color_data = 12'b011001111001;
		if(({row_reg, col_reg}==18'b000111101001100110)) color_data = 12'b011110001000;
		if(({row_reg, col_reg}==18'b000111101001100111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b000111101001101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b000111101001101001) && ({row_reg, col_reg}<18'b000111101001110110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b000111101001110110) && ({row_reg, col_reg}<18'b000111101001111001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b000111101001111001)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b000111101001111010) && ({row_reg, col_reg}<18'b000111101001111100)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}>=18'b000111101001111100) && ({row_reg, col_reg}<18'b000111101010000100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b000111101010000100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b000111101010000101) && ({row_reg, col_reg}<18'b000111101010000111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b000111101010000111)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b000111101010001000) && ({row_reg, col_reg}<18'b000111101010001010)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b000111101010001010)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b000111101010001011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b000111101010001100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b000111101010001101)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b000111101010001110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b000111101010001111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b000111101010010000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b000111101010010001)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b000111101010010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b000111101010010011) && ({row_reg, col_reg}<18'b000111101010010110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b000111101010010110)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b000111101010010111)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}>=18'b000111101010011000) && ({row_reg, col_reg}<18'b000111101010011011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b000111101010011011)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b000111101010011100) && ({row_reg, col_reg}<18'b000111101010100000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b000111101010100000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b000111101010100001)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}==18'b000111101010100010)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==18'b000111101010100011)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b000111101010100100)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}==18'b000111101010100101)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b000111101010100110)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}>=18'b000111101010100111) && ({row_reg, col_reg}<18'b000111101010101001)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b000111101010101001) && ({row_reg, col_reg}<18'b000111101010101100)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b000111101010101100) && ({row_reg, col_reg}<18'b000111110001011100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b000111110001011100) && ({row_reg, col_reg}<18'b000111110001100000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b000111110001100000) && ({row_reg, col_reg}<18'b000111110001100010)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b000111110001100010)) color_data = 12'b011110011011;
		if(({row_reg, col_reg}==18'b000111110001100011)) color_data = 12'b011010001001;
		if(({row_reg, col_reg}==18'b000111110001100100)) color_data = 12'b011110001001;
		if(({row_reg, col_reg}==18'b000111110001100101)) color_data = 12'b011110001000;
		if(({row_reg, col_reg}==18'b000111110001100110)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==18'b000111110001100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b000111110001101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b000111110001101001)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}>=18'b000111110001101010) && ({row_reg, col_reg}<18'b000111110001110000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b000111110001110000) && ({row_reg, col_reg}<18'b000111110001110100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b000111110001110100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b000111110001110101) && ({row_reg, col_reg}<18'b000111110001111010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b000111110001111010) && ({row_reg, col_reg}<18'b000111110010000100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b000111110010000100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b000111110010000101) && ({row_reg, col_reg}<18'b000111110010001001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b000111110010001001)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b000111110010001010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b000111110010001011) && ({row_reg, col_reg}<18'b000111110010001101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b000111110010001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b000111110010001110) && ({row_reg, col_reg}<18'b000111110010010000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b000111110010010000) && ({row_reg, col_reg}<18'b000111110010010011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b000111110010010011)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b000111110010010100) && ({row_reg, col_reg}<18'b000111110010010110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b000111110010010110)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b000111110010010111)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b000111110010011000) && ({row_reg, col_reg}<18'b000111110010011100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b000111110010011100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b000111110010011101) && ({row_reg, col_reg}<18'b000111110010100000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b000111110010100000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b000111110010100001) && ({row_reg, col_reg}<18'b000111110010100100)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}==18'b000111110010100100)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}>=18'b000111110010100101) && ({row_reg, col_reg}<18'b000111110010100111)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b000111110010100111)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}>=18'b000111110010101000) && ({row_reg, col_reg}<18'b000111110010101010)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b000111110010101010) && ({row_reg, col_reg}<18'b000111110010101110)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b000111110010101110) && ({row_reg, col_reg}<18'b000111111001011001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b000111111001011001) && ({row_reg, col_reg}<18'b000111111001100000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b000111111001100000) && ({row_reg, col_reg}<18'b000111111001100010)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b000111111001100010)) color_data = 12'b100010011011;
		if(({row_reg, col_reg}==18'b000111111001100011)) color_data = 12'b011001111001;
		if(({row_reg, col_reg}==18'b000111111001100100)) color_data = 12'b011110001001;
		if(({row_reg, col_reg}==18'b000111111001100101)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==18'b000111111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b000111111001100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b000111111001101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b000111111001101001)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b000111111001101010) && ({row_reg, col_reg}<18'b000111111001101100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b000111111001101100) && ({row_reg, col_reg}<18'b000111111001101111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b000111111001101111) && ({row_reg, col_reg}<18'b000111111001111010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b000111111001111010) && ({row_reg, col_reg}<18'b000111111001111111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b000111111001111111)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}>=18'b000111111010000000) && ({row_reg, col_reg}<18'b000111111010000100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b000111111010000100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b000111111010000101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b000111111010000110) && ({row_reg, col_reg}<18'b000111111010001000)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b000111111010001000) && ({row_reg, col_reg}<18'b000111111010001101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b000111111010001101)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b000111111010001110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b000111111010001111) && ({row_reg, col_reg}<18'b000111111010010011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b000111111010010011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b000111111010010100) && ({row_reg, col_reg}<18'b000111111010010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b000111111010010110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b000111111010010111)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b000111111010011000) && ({row_reg, col_reg}<18'b000111111010011011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b000111111010011011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b000111111010011100) && ({row_reg, col_reg}<18'b000111111010100000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b000111111010100000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b000111111010100001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b000111111010100010)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}==18'b000111111010100011)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}>=18'b000111111010100100) && ({row_reg, col_reg}<18'b000111111010100110)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b000111111010100110)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}==18'b000111111010100111)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b000111111010101000)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}==18'b000111111010101001)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b000111111010101010) && ({row_reg, col_reg}<18'b000111111010101110)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b000111111010101110) && ({row_reg, col_reg}<18'b001000000001010000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001000000001010000)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}==18'b001000000001010001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001000000001010010) && ({row_reg, col_reg}<18'b001000000001010100)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001000000001010100) && ({row_reg, col_reg}<18'b001000000001011001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001000000001011001)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001000000001011010) && ({row_reg, col_reg}<18'b001000000001011100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001000000001011100)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001000000001011101)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001000000001011110)) color_data = 12'b011110011100;
		if(({row_reg, col_reg}==18'b001000000001011111)) color_data = 12'b011110011011;
		if(({row_reg, col_reg}>=18'b001000000001100000) && ({row_reg, col_reg}<18'b001000000001100010)) color_data = 12'b100010011010;
		if(({row_reg, col_reg}>=18'b001000000001100010) && ({row_reg, col_reg}<18'b001000000001100100)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}==18'b001000000001100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b001000000001100101) && ({row_reg, col_reg}<18'b001000000001100111)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b001000000001100111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001000000001101000) && ({row_reg, col_reg}<18'b001000000001101110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b001000000001101110) && ({row_reg, col_reg}<18'b001000000001110001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001000000001110001) && ({row_reg, col_reg}<18'b001000000001111111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001000000001111111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001000000010000000) && ({row_reg, col_reg}<18'b001000000010000010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b001000000010000010)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001000000010000011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b001000000010000100) && ({row_reg, col_reg}<18'b001000000010000110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001000000010000110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001000000010000111) && ({row_reg, col_reg}<18'b001000000010001001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001000000010001001)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b001000000010001010) && ({row_reg, col_reg}<18'b001000000010001100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001000000010001100)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001000000010001101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b001000000010001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b001000000010001111) && ({row_reg, col_reg}<18'b001000000010010010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001000000010010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b001000000010010011) && ({row_reg, col_reg}<18'b001000000010010110)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b001000000010010110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b001000000010010111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001000000010011000) && ({row_reg, col_reg}<18'b001000000010011100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001000000010011100) && ({row_reg, col_reg}<18'b001000000010011110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001000000010011110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001000000010011111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b001000000010100000) && ({row_reg, col_reg}<18'b001000000010100011)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001000000010100011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b001000000010100100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001000000010100101)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}==18'b001000000010100110)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=18'b001000000010100111) && ({row_reg, col_reg}<18'b001000000010101001)) color_data = 12'b100010011010;
		if(({row_reg, col_reg}==18'b001000000010101001)) color_data = 12'b011110011011;
		if(({row_reg, col_reg}==18'b001000000010101010)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b001000000010101011)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b001000000010101100) && ({row_reg, col_reg}<18'b001000000010110101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001000000010110101) && ({row_reg, col_reg}<18'b001000000010111000)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b001000000010111000) && ({row_reg, col_reg}<18'b001000001001010010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001000001001010010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001000001001010011) && ({row_reg, col_reg}<18'b001000001001011001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001000001001011001)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001000001001011010) && ({row_reg, col_reg}<18'b001000001001011101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001000001001011101)) color_data = 12'b011110011101;
		if(({row_reg, col_reg}==18'b001000001001011110)) color_data = 12'b011010001011;
		if(({row_reg, col_reg}==18'b001000001001011111)) color_data = 12'b011010001010;
		if(({row_reg, col_reg}==18'b001000001001100000)) color_data = 12'b011110001000;
		if(({row_reg, col_reg}==18'b001000001001100001)) color_data = 12'b011110001001;
		if(({row_reg, col_reg}==18'b001000001001100010)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=18'b001000001001100011) && ({row_reg, col_reg}<18'b001000001001100111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001000001001100111) && ({row_reg, col_reg}<18'b001000001001111011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b001000001001111011) && ({row_reg, col_reg}<18'b001000001001111111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001000001001111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b001000001010000000) && ({row_reg, col_reg}<18'b001000001010000011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001000001010000011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001000001010000100)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b001000001010000101) && ({row_reg, col_reg}<18'b001000001010001000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001000001010001000) && ({row_reg, col_reg}<18'b001000001010001010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001000001010001010)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001000001010001011) && ({row_reg, col_reg}<18'b001000001010001101)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b001000001010001101) && ({row_reg, col_reg}<18'b001000001010010000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001000001010010000) && ({row_reg, col_reg}<18'b001000001010010010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b001000001010010010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001000001010010011) && ({row_reg, col_reg}<18'b001000001010010101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001000001010010101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001000001010010110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001000001010010111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001000001010011000) && ({row_reg, col_reg}<18'b001000001010011010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b001000001010011010) && ({row_reg, col_reg}<18'b001000001010011100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001000001010011100) && ({row_reg, col_reg}<18'b001000001010011110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001000001010011110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001000001010011111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b001000001010100000) && ({row_reg, col_reg}<18'b001000001010100011)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001000001010100011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b001000001010100100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001000001010100101)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}==18'b001000001010100110)) color_data = 12'b011110001000;
		if(({row_reg, col_reg}>=18'b001000001010100111) && ({row_reg, col_reg}<18'b001000001010101001)) color_data = 12'b011110001001;
		if(({row_reg, col_reg}==18'b001000001010101001)) color_data = 12'b011010001010;
		if(({row_reg, col_reg}==18'b001000001010101010)) color_data = 12'b011110011100;
		if(({row_reg, col_reg}==18'b001000001010101011)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b001000001010101100) && ({row_reg, col_reg}<18'b001000001010110101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001000001010110101) && ({row_reg, col_reg}<18'b001000001010111000)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b001000001010111000) && ({row_reg, col_reg}<18'b001000010001010100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001000010001010100)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b001000010001010101) && ({row_reg, col_reg}<18'b001000010001011011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001000010001011011) && ({row_reg, col_reg}<18'b001000010001011101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001000010001011101)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001000010001011110)) color_data = 12'b011010001011;
		if(({row_reg, col_reg}==18'b001000010001011111)) color_data = 12'b011001111001;
		if(({row_reg, col_reg}==18'b001000010001100000)) color_data = 12'b011001111000;
		if(({row_reg, col_reg}==18'b001000010001100001)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==18'b001000010001100010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b001000010001100011)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b001000010001100100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001000010001100101) && ({row_reg, col_reg}<18'b001000010001111011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b001000010001111011) && ({row_reg, col_reg}<18'b001000010001111101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001000010001111101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001000010001111110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001000010001111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b001000010010000000) && ({row_reg, col_reg}<18'b001000010010000100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001000010010000100)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b001000010010000101) && ({row_reg, col_reg}<18'b001000010010000111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001000010010000111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001000010010001000)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b001000010010001001) && ({row_reg, col_reg}<18'b001000010010001110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001000010010001110)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001000010010001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001000010010010000) && ({row_reg, col_reg}<18'b001000010010010010)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001000010010010010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001000010010010011) && ({row_reg, col_reg}<18'b001000010010011001)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b001000010010011001) && ({row_reg, col_reg}<18'b001000010010011100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001000010010011100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b001000010010011101) && ({row_reg, col_reg}<18'b001000010010011111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001000010010011111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001000010010100000)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001000010010100001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001000010010100010)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001000010010100011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001000010010100100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001000010010100101)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}==18'b001000010010100110)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==18'b001000010010100111)) color_data = 12'b011110001000;
		if(({row_reg, col_reg}==18'b001000010010101000)) color_data = 12'b011001111000;
		if(({row_reg, col_reg}==18'b001000010010101001)) color_data = 12'b011010001001;
		if(({row_reg, col_reg}==18'b001000010010101010)) color_data = 12'b011110011011;
		if(({row_reg, col_reg}==18'b001000010010101011)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b001000010010101100) && ({row_reg, col_reg}<18'b001000010010101111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001000010010101111)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b001000010010110000) && ({row_reg, col_reg}<18'b001000010010110101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001000010010110101) && ({row_reg, col_reg}<18'b001000010010111000)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b001000010010111000) && ({row_reg, col_reg}<18'b001000011001011011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001000011001011011) && ({row_reg, col_reg}<18'b001000011001011101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001000011001011101)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}==18'b001000011001011110)) color_data = 12'b011010001011;
		if(({row_reg, col_reg}==18'b001000011001011111)) color_data = 12'b011001111001;
		if(({row_reg, col_reg}==18'b001000011001100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001000011001100001)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==18'b001000011001100010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b001000011001100011)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}>=18'b001000011001100100) && ({row_reg, col_reg}<18'b001000011001100111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001000011001100111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b001000011001101000) && ({row_reg, col_reg}<18'b001000011001101010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001000011001101010) && ({row_reg, col_reg}<18'b001000011001111011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001000011001111011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001000011001111100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001000011001111101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001000011001111110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001000011001111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b001000011010000000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001000011010000001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b001000011010000010) && ({row_reg, col_reg}<18'b001000011010000100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001000011010000100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b001000011010000101) && ({row_reg, col_reg}<18'b001000011010000111)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001000011010000111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001000011010001000) && ({row_reg, col_reg}<18'b001000011010010000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001000011010010000)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001000011010010001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001000011010010010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001000011010010011) && ({row_reg, col_reg}<18'b001000011010011010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b001000011010011010) && ({row_reg, col_reg}<18'b001000011010011101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001000011010011101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001000011010011110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001000011010011111) && ({row_reg, col_reg}<18'b001000011010100001)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001000011010100001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001000011010100010)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}>=18'b001000011010100011) && ({row_reg, col_reg}<18'b001000011010100101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001000011010100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b001000011010100110) && ({row_reg, col_reg}<18'b001000011010101000)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==18'b001000011010101000)) color_data = 12'b011110001000;
		if(({row_reg, col_reg}==18'b001000011010101001)) color_data = 12'b011110001001;
		if(({row_reg, col_reg}==18'b001000011010101010)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}==18'b001000011010101011)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001000011010101100)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001000011010101101) && ({row_reg, col_reg}<18'b001000011010110001)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b001000011010110001) && ({row_reg, col_reg}<18'b001000011010110101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001000011010110101) && ({row_reg, col_reg}<18'b001000011010110111)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b001000011010110111) && ({row_reg, col_reg}<18'b001000100001010000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001000100001010000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001000100001010001) && ({row_reg, col_reg}<18'b001000100001011000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001000100001011000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001000100001011001) && ({row_reg, col_reg}<18'b001000100001011011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001000100001011011)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001000100001011100)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001000100001011101)) color_data = 12'b011110011100;
		if(({row_reg, col_reg}==18'b001000100001011110)) color_data = 12'b011110001010;
		if(({row_reg, col_reg}==18'b001000100001011111)) color_data = 12'b011110001001;
		if(({row_reg, col_reg}==18'b001000100001100000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b001000100001100001) && ({row_reg, col_reg}<18'b001000100001100011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b001000100001100011) && ({row_reg, col_reg}<18'b001000100001101001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001000100001101001) && ({row_reg, col_reg}<18'b001000100001111010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001000100001111010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001000100001111011) && ({row_reg, col_reg}<18'b001000100001111110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001000100001111110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b001000100001111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b001000100010000000) && ({row_reg, col_reg}<18'b001000100010000100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001000100010000100)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}>=18'b001000100010000101) && ({row_reg, col_reg}<18'b001000100010000111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001000100010000111)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001000100010001000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001000100010001001)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b001000100010001010) && ({row_reg, col_reg}<18'b001000100010001100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001000100010001100)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b001000100010001101) && ({row_reg, col_reg}<18'b001000100010010000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001000100010010000)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b001000100010010001) && ({row_reg, col_reg}<18'b001000100010010011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001000100010010011) && ({row_reg, col_reg}<18'b001000100010011100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001000100010011100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001000100010011101) && ({row_reg, col_reg}<18'b001000100010100001)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001000100010100001)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b001000100010100010) && ({row_reg, col_reg}<18'b001000100010100101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001000100010100101) && ({row_reg, col_reg}<18'b001000100010100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b001000100010100111) && ({row_reg, col_reg}<18'b001000100010101001)) color_data = 12'b011110001000;
		if(({row_reg, col_reg}==18'b001000100010101001)) color_data = 12'b011010001001;
		if(({row_reg, col_reg}==18'b001000100010101010)) color_data = 12'b011110011011;
		if(({row_reg, col_reg}==18'b001000100010101011)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001000100010101100)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001000100010101101) && ({row_reg, col_reg}<18'b001000100010110010)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b001000100010110010) && ({row_reg, col_reg}<18'b001000100010110101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001000100010110101) && ({row_reg, col_reg}<18'b001000100010110111)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b001000100010110111) && ({row_reg, col_reg}<18'b001000101001010000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001000101001010000) && ({row_reg, col_reg}<18'b001000101001010010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001000101001010010) && ({row_reg, col_reg}<18'b001000101001010111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001000101001010111) && ({row_reg, col_reg}<18'b001000101001011100)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001000101001011100)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001000101001011101)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b001000101001011110)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}==18'b001000101001011111)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}>=18'b001000101001100000) && ({row_reg, col_reg}<18'b001000101001100011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001000101001100011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001000101001100100) && ({row_reg, col_reg}<18'b001000101001100110)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}>=18'b001000101001100110) && ({row_reg, col_reg}<18'b001000101001101001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001000101001101001) && ({row_reg, col_reg}<18'b001000101001110101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b001000101001110101) && ({row_reg, col_reg}<18'b001000101001110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001000101001110111)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001000101001111000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001000101001111001) && ({row_reg, col_reg}<18'b001000101001111011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001000101001111011)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b001000101001111100) && ({row_reg, col_reg}<18'b001000101001111111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001000101001111111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001000101010000000) && ({row_reg, col_reg}<18'b001000101010000100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001000101010000100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b001000101010000101) && ({row_reg, col_reg}<18'b001000101010001001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001000101010001001) && ({row_reg, col_reg}<18'b001000101010001011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b001000101010001011) && ({row_reg, col_reg}<18'b001000101010001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001000101010001111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001000101010010000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001000101010010001) && ({row_reg, col_reg}<18'b001000101010011100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001000101010011100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001000101010011101) && ({row_reg, col_reg}<18'b001000101010100000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001000101010100000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001000101010100001) && ({row_reg, col_reg}<18'b001000101010100101)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b001000101010100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b001000101010100110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001000101010100111)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b001000101010101000)) color_data = 12'b011110001000;
		if(({row_reg, col_reg}==18'b001000101010101001)) color_data = 12'b011110001001;
		if(({row_reg, col_reg}==18'b001000101010101010)) color_data = 12'b011110011011;
		if(({row_reg, col_reg}==18'b001000101010101011)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}>=18'b001000101010101100) && ({row_reg, col_reg}<18'b001000101010101110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001000101010101110) && ({row_reg, col_reg}<18'b001000101010110010)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b001000101010110010) && ({row_reg, col_reg}<18'b001000101010110101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001000101010110101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001000101010110110)) color_data = 12'b011010101101;

		if(({row_reg, col_reg}>=18'b001000101010110111) && ({row_reg, col_reg}<18'b001000110001010000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001000110001010000) && ({row_reg, col_reg}<18'b001000110001010010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001000110001010010) && ({row_reg, col_reg}<18'b001000110001011010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001000110001011010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001000110001011011)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001000110001011100)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}==18'b001000110001011101)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b001000110001011110)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b001000110001011111)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}>=18'b001000110001100000) && ({row_reg, col_reg}<18'b001000110001100100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b001000110001100100) && ({row_reg, col_reg}<18'b001000110001101001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001000110001101001) && ({row_reg, col_reg}<18'b001000110001110101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001000110001110101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001000110001110110) && ({row_reg, col_reg}<18'b001000110001111010)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001000110001111010)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b001000110001111011) && ({row_reg, col_reg}<18'b001000110010000011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001000110010000011)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b001000110010000100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001000110010000101)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001000110010000110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001000110010000111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001000110010001000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001000110010001001) && ({row_reg, col_reg}<18'b001000110010011100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001000110010011100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001000110010011101) && ({row_reg, col_reg}<18'b001000110010100000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001000110010100000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001000110010100001) && ({row_reg, col_reg}<18'b001000110010100111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001000110010100111)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b001000110010101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001000110010101001)) color_data = 12'b011110001001;
		if(({row_reg, col_reg}==18'b001000110010101010)) color_data = 12'b100010011011;
		if(({row_reg, col_reg}==18'b001000110010101011)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b001000110010101100)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b001000110010101101) && ({row_reg, col_reg}<18'b001000110010101111)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001000110010101111) && ({row_reg, col_reg}<18'b001000110010110001)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b001000110010110001) && ({row_reg, col_reg}<18'b001000110010110101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001000110010110101) && ({row_reg, col_reg}<18'b001000110010111000)) color_data = 12'b011010101101;

		if(({row_reg, col_reg}>=18'b001000110010111000) && ({row_reg, col_reg}<18'b001000111001010000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001000111001010000) && ({row_reg, col_reg}<18'b001000111001010010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001000111001010010) && ({row_reg, col_reg}<18'b001000111001011000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001000111001011000) && ({row_reg, col_reg}<18'b001000111001011010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001000111001011010) && ({row_reg, col_reg}<18'b001000111001011100)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001000111001011100)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}==18'b001000111001011101)) color_data = 12'b100010011011;
		if(({row_reg, col_reg}==18'b001000111001011110)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b001000111001011111)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}>=18'b001000111001100000) && ({row_reg, col_reg}<18'b001000111001100101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b001000111001100101) && ({row_reg, col_reg}<18'b001000111001101001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001000111001101001) && ({row_reg, col_reg}<18'b001000111001110101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001000111001110101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001000111001110110) && ({row_reg, col_reg}<18'b001000111001111000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001000111001111000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001000111001111001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001000111001111010)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b001000111001111011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b001000111001111100) && ({row_reg, col_reg}<18'b001000111010000100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001000111010000100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b001000111010000101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001000111010000110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001000111010000111)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001000111010001000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001000111010001001) && ({row_reg, col_reg}<18'b001000111010011100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001000111010011100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001000111010011101) && ({row_reg, col_reg}<18'b001000111010100000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001000111010100000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001000111010100001) && ({row_reg, col_reg}<18'b001000111010100111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b001000111010100111) && ({row_reg, col_reg}<18'b001000111010101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001000111010101001)) color_data = 12'b011110001000;
		if(({row_reg, col_reg}==18'b001000111010101010)) color_data = 12'b100010011010;
		if(({row_reg, col_reg}==18'b001000111010101011)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}==18'b001000111010101100)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}==18'b001000111010101101)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001000111010101110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001000111010101111) && ({row_reg, col_reg}<18'b001000111010110101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001000111010110101) && ({row_reg, col_reg}<18'b001000111010110111)) color_data = 12'b011010101101;

		if(({row_reg, col_reg}>=18'b001000111010110111) && ({row_reg, col_reg}<18'b001001000001010000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001001000001010000) && ({row_reg, col_reg}<18'b001001000001010010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001001000001010010) && ({row_reg, col_reg}<18'b001001000001010111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001001000001010111) && ({row_reg, col_reg}<18'b001001000001011001)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001001000001011001) && ({row_reg, col_reg}<18'b001001000001011011)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001001000001011011)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}==18'b001001000001011100)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b001001000001011101)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}>=18'b001001000001011110) && ({row_reg, col_reg}<18'b001001000001100000)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}>=18'b001001000001100000) && ({row_reg, col_reg}<18'b001001000001100010)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}>=18'b001001000001100010) && ({row_reg, col_reg}<18'b001001000001100100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b001001000001100100) && ({row_reg, col_reg}<18'b001001000001101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001001000001101000) && ({row_reg, col_reg}<18'b001001000001110110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001001000001110110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001001000001110111) && ({row_reg, col_reg}<18'b001001000001111001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001001000001111001)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001001000001111010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b001001000001111011) && ({row_reg, col_reg}<18'b001001000010000010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001001000010000010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b001001000010000011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001001000010000100)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b001001000010000101) && ({row_reg, col_reg}<18'b001001000010001001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001001000010001001)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001001000010001010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001001000010001011) && ({row_reg, col_reg}<18'b001001000010011100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001001000010011100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001001000010011101) && ({row_reg, col_reg}<18'b001001000010100000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001001000010100000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001001000010100001) && ({row_reg, col_reg}<18'b001001000010101000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001001000010101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001001000010101001)) color_data = 12'b011110001000;
		if(({row_reg, col_reg}==18'b001001000010101010)) color_data = 12'b100010011010;
		if(({row_reg, col_reg}==18'b001001000010101011)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b001001000010101100)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}>=18'b001001000010101101) && ({row_reg, col_reg}<18'b001001000010101111)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b001001000010101111) && ({row_reg, col_reg}<18'b001001000010110010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001001000010110010) && ({row_reg, col_reg}<18'b001001000010110100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001001000010110100)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b001001000010110101) && ({row_reg, col_reg}<18'b001001001001010000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001001001001010000) && ({row_reg, col_reg}<18'b001001001001010010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001001001001010010) && ({row_reg, col_reg}<18'b001001001001010110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001001001001010110) && ({row_reg, col_reg}<18'b001001001001011001)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001001001001011001)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001001001001011010)) color_data = 12'b011110011100;
		if(({row_reg, col_reg}==18'b001001001001011011)) color_data = 12'b011110011011;
		if(({row_reg, col_reg}==18'b001001001001011100)) color_data = 12'b100010011011;
		if(({row_reg, col_reg}==18'b001001001001011101)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}==18'b001001001001011110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001001001001011111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==18'b001001001001100000)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}>=18'b001001001001100001) && ({row_reg, col_reg}<18'b001001001001110000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001001001001110000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001001001001110001) && ({row_reg, col_reg}<18'b001001001001110101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001001001001110101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001001001001110110) && ({row_reg, col_reg}<18'b001001001001111000)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b001001001001111000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b001001001001111001)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b001001001001111010)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b001001001001111011) && ({row_reg, col_reg}<18'b001001001001111111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001001001001111111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001001001010000000) && ({row_reg, col_reg}<18'b001001001010000100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b001001001010000100) && ({row_reg, col_reg}<18'b001001001010000111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001001001010000111) && ({row_reg, col_reg}<18'b001001001010001001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001001001010001001) && ({row_reg, col_reg}<18'b001001001010011110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001001001010011110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001001001010011111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001001001010100000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001001001010100001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001001001010100010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001001001010100011) && ({row_reg, col_reg}<18'b001001001010100111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b001001001010100111) && ({row_reg, col_reg}<18'b001001001010101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b001001001010101001)) color_data = 12'b011110001000;
		if(({row_reg, col_reg}==18'b001001001010101010)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}==18'b001001001010101011)) color_data = 12'b100010011010;
		if(({row_reg, col_reg}>=18'b001001001010101100) && ({row_reg, col_reg}<18'b001001001010101110)) color_data = 12'b011110011011;
		if(({row_reg, col_reg}==18'b001001001010101110)) color_data = 12'b011110011100;
		if(({row_reg, col_reg}==18'b001001001010101111)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b001001001010110000) && ({row_reg, col_reg}<18'b001001001010110100)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b001001001010110100) && ({row_reg, col_reg}<18'b001001010001010000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001001010001010000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001001010001010001) && ({row_reg, col_reg}<18'b001001010001010110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001001010001010110) && ({row_reg, col_reg}<18'b001001010001011000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001001010001011000)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001001010001011001)) color_data = 12'b011010011011;
		if(({row_reg, col_reg}==18'b001001010001011010)) color_data = 12'b011010001010;
		if(({row_reg, col_reg}==18'b001001010001011011)) color_data = 12'b011010001001;
		if(({row_reg, col_reg}==18'b001001010001011100)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==18'b001001010001011101)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}==18'b001001010001011110)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}==18'b001001010001011111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001001010001100000)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}>=18'b001001010001100001) && ({row_reg, col_reg}<18'b001001010001101110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b001001010001101110) && ({row_reg, col_reg}<18'b001001010001110000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001001010001110000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001001010001110001)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b001001010001110010) && ({row_reg, col_reg}<18'b001001010001110101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001001010001110101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b001001010001110110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001001010001110111) && ({row_reg, col_reg}<18'b001001010001111001)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001001010001111001)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b001001010001111010) && ({row_reg, col_reg}<18'b001001010001111110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001001010001111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001001010001111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b001001010010000000) && ({row_reg, col_reg}<18'b001001010010000011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001001010010000011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b001001010010000100) && ({row_reg, col_reg}<18'b001001010010011110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001001010010011110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001001010010011111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001001010010100000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001001010010100001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001001010010100010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001001010010100011) && ({row_reg, col_reg}<18'b001001010010100111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001001010010100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b001001010010101000) && ({row_reg, col_reg}<18'b001001010010101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001001010010101010)) color_data = 12'b011110001000;
		if(({row_reg, col_reg}==18'b001001010010101011)) color_data = 12'b011110001001;
		if(({row_reg, col_reg}==18'b001001010010101100)) color_data = 12'b011001111001;
		if(({row_reg, col_reg}==18'b001001010010101101)) color_data = 12'b011010001001;
		if(({row_reg, col_reg}==18'b001001010010101110)) color_data = 12'b011010001010;
		if(({row_reg, col_reg}==18'b001001010010101111)) color_data = 12'b011110011100;
		if(({row_reg, col_reg}>=18'b001001010010110000) && ({row_reg, col_reg}<18'b001001010010110101)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b001001010010110101) && ({row_reg, col_reg}<18'b001001011001010000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001001011001010000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001001011001010001) && ({row_reg, col_reg}<18'b001001011001010110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001001011001010110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001001011001010111) && ({row_reg, col_reg}<18'b001001011001011001)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001001011001011001)) color_data = 12'b011010001011;
		if(({row_reg, col_reg}==18'b001001011001011010)) color_data = 12'b011010001001;
		if(({row_reg, col_reg}==18'b001001011001011011)) color_data = 12'b011110001001;
		if(({row_reg, col_reg}==18'b001001011001011100)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==18'b001001011001011101)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}==18'b001001011001011110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001001011001011111) && ({row_reg, col_reg}<18'b001001011001101110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b001001011001101110) && ({row_reg, col_reg}<18'b001001011001110000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001001011001110000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b001001011001110001) && ({row_reg, col_reg}<18'b001001011001110101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001001011001110101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b001001011001110110) && ({row_reg, col_reg}<18'b001001011001111110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001001011001111110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b001001011001111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b001001011010000000)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001001011010000001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001001011010000010) && ({row_reg, col_reg}<18'b001001011010000100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001001011010000100) && ({row_reg, col_reg}<18'b001001011010011010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001001011010011010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001001011010011011) && ({row_reg, col_reg}<18'b001001011010011110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001001011010011110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001001011010011111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001001011010100000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001001011010100001) && ({row_reg, col_reg}<18'b001001011010101000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b001001011010101000) && ({row_reg, col_reg}<18'b001001011010101101)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==18'b001001011010101101)) color_data = 12'b011110001001;
		if(({row_reg, col_reg}==18'b001001011010101110)) color_data = 12'b011010001001;
		if(({row_reg, col_reg}==18'b001001011010101111)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b001001011010110000)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b001001011010110001) && ({row_reg, col_reg}<18'b001001011010110101)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b001001011010110101) && ({row_reg, col_reg}<18'b001001100001010101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001001100001010101) && ({row_reg, col_reg}<18'b001001100001011000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001001100001011000)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}==18'b001001100001011001)) color_data = 12'b011010001010;
		if(({row_reg, col_reg}==18'b001001100001011010)) color_data = 12'b011001111001;
		if(({row_reg, col_reg}>=18'b001001100001011011) && ({row_reg, col_reg}<18'b001001100001011101)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==18'b001001100001011101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b001001100001011110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001001100001011111) && ({row_reg, col_reg}<18'b001001100001101100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001001100001101100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001001100001101101) && ({row_reg, col_reg}<18'b001001100001101111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001001100001101111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001001100001110000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001001100001110001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001001100001110010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001001100001110011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b001001100001110100) && ({row_reg, col_reg}<18'b001001100001110110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001001100001110110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001001100001110111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b001001100001111000) && ({row_reg, col_reg}<18'b001001100001111111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001001100001111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b001001100010000000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001001100010000001)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b001001100010000010) && ({row_reg, col_reg}<18'b001001100010000100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001001100010000100) && ({row_reg, col_reg}<18'b001001100010010000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b001001100010010000) && ({row_reg, col_reg}<18'b001001100010010010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001001100010010010) && ({row_reg, col_reg}<18'b001001100010011101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001001100010011101)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==18'b001001100010011110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001001100010011111)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==18'b001001100010100000)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001001100010100001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001001100010100010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001001100010100011) && ({row_reg, col_reg}<18'b001001100010101001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001001100010101001)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==18'b001001100010101010)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}>=18'b001001100010101011) && ({row_reg, col_reg}<18'b001001100010101101)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==18'b001001100010101101)) color_data = 12'b011110001001;
		if(({row_reg, col_reg}==18'b001001100010101110)) color_data = 12'b011010001001;
		if(({row_reg, col_reg}==18'b001001100010101111)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b001001100010110000)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b001001100010110001) && ({row_reg, col_reg}<18'b001001100010110101)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b001001100010110101) && ({row_reg, col_reg}<18'b001001101001010101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001001101001010101) && ({row_reg, col_reg}<18'b001001101001010111)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001001101001010111)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001001101001011000)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}==18'b001001101001011001)) color_data = 12'b011110011010;
		if(({row_reg, col_reg}==18'b001001101001011010)) color_data = 12'b011001111001;
		if(({row_reg, col_reg}==18'b001001101001011011)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==18'b001001101001011100)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}==18'b001001101001011101)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b001001101001011110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001001101001011111) && ({row_reg, col_reg}<18'b001001101001101100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001001101001101100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001001101001101101) && ({row_reg, col_reg}<18'b001001101001110001)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b001001101001110001) && ({row_reg, col_reg}<18'b001001101001110101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001001101001110101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b001001101001110110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b001001101001110111) && ({row_reg, col_reg}<18'b001001101001111001)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001001101001111001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b001001101001111010) && ({row_reg, col_reg}<18'b001001101001111100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001001101001111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001001101001111101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001001101001111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001001101001111111)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b001001101010000000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001001101010000001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001001101010000010) && ({row_reg, col_reg}<18'b001001101010000100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001001101010000100) && ({row_reg, col_reg}<18'b001001101010011100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001001101010011100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001001101010011101) && ({row_reg, col_reg}<18'b001001101010100000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001001101010100000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001001101010100001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001001101010100010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001001101010100011) && ({row_reg, col_reg}<18'b001001101010101100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001001101010101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001001101010101101)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==18'b001001101010101110)) color_data = 12'b011010001001;
		if(({row_reg, col_reg}==18'b001001101010101111)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b001001101010110000)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b001001101010110001) && ({row_reg, col_reg}<18'b001001101010110100)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b001001101010110100) && ({row_reg, col_reg}<18'b001001110001010101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001001110001010101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001001110001010110) && ({row_reg, col_reg}<18'b001001110001011000)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001001110001011000)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b001001110001011001)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}==18'b001001110001011010)) color_data = 12'b100010011010;
		if(({row_reg, col_reg}==18'b001001110001011011)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}==18'b001001110001011100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b001001110001011101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001001110001011110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001001110001011111) && ({row_reg, col_reg}<18'b001001110001101100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b001001110001101100) && ({row_reg, col_reg}<18'b001001110001110001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001001110001110001)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b001001110001110010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001001110001110011)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b001001110001110100) && ({row_reg, col_reg}<18'b001001110001110110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b001001110001110110) && ({row_reg, col_reg}<18'b001001110001111010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001001110001111010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b001001110001111011) && ({row_reg, col_reg}<18'b001001110001111111)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b001001110001111111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b001001110010000000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001001110010000001)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b001001110010000010) && ({row_reg, col_reg}<18'b001001110010000100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001001110010000100) && ({row_reg, col_reg}<18'b001001110010011011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001001110010011011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001001110010011100) && ({row_reg, col_reg}<18'b001001110010011110)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==18'b001001110010011110)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b001001110010011111)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==18'b001001110010100000)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b001001110010100001) && ({row_reg, col_reg}<18'b001001110010101100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001001110010101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001001110010101101)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==18'b001001110010101110)) color_data = 12'b011110001001;
		if(({row_reg, col_reg}==18'b001001110010101111)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}==18'b001001110010110000)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b001001110010110001) && ({row_reg, col_reg}<18'b001001110010110100)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001001110010110100) && ({row_reg, col_reg}<18'b001001110010110110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001001110010110110)) color_data = 12'b011010101111;

		if(({row_reg, col_reg}>=18'b001001110010110111) && ({row_reg, col_reg}<18'b001001111001010011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001001111001010011)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}>=18'b001001111001010100) && ({row_reg, col_reg}<18'b001001111001010110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001001111001010110) && ({row_reg, col_reg}<18'b001001111001011000)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001001111001011000)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b001001111001011001)) color_data = 12'b100110111100;
		if(({row_reg, col_reg}==18'b001001111001011010)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b001001111001011011)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}>=18'b001001111001011100) && ({row_reg, col_reg}<18'b001001111001011111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001001111001011111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001001111001100000) && ({row_reg, col_reg}<18'b001001111001101000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b001001111001101000) && ({row_reg, col_reg}<18'b001001111001101011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001001111001101011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b001001111001101100) && ({row_reg, col_reg}<18'b001001111001110001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001001111001110001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001001111001110010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b001001111001110011) && ({row_reg, col_reg}<18'b001001111001110110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001001111001110110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b001001111001110111) && ({row_reg, col_reg}<18'b001001111001111010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001001111001111010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001001111001111011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001001111001111100) && ({row_reg, col_reg}<18'b001001111010000000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001001111010000000) && ({row_reg, col_reg}<18'b001001111010000010)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b001001111010000010) && ({row_reg, col_reg}<18'b001001111010000100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001001111010000100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001001111010000101) && ({row_reg, col_reg}<18'b001001111010011001)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001001111010011001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001001111010011010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001001111010011011)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001001111010011100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b001001111010011101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001001111010011110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001001111010011111) && ({row_reg, col_reg}<18'b001001111010100010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001001111010100010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b001001111010100011) && ({row_reg, col_reg}<18'b001001111010101101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001001111010101101)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==18'b001001111010101110)) color_data = 12'b011101111001;
		if(({row_reg, col_reg}==18'b001001111010101111)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}>=18'b001001111010110000) && ({row_reg, col_reg}<18'b001001111010110100)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001001111010110100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001001111010110101)) color_data = 12'b011010101111;

		if(({row_reg, col_reg}>=18'b001001111010110110) && ({row_reg, col_reg}<18'b001010000001010010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001010000001010010) && ({row_reg, col_reg}<18'b001010000001010100)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b001010000001010100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001010000001010101) && ({row_reg, col_reg}<18'b001010000001010111)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001010000001010111)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001010000001011000)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b001010000001011001)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==18'b001010000001011010)) color_data = 12'b101010111011;
		if(({row_reg, col_reg}==18'b001010000001011011)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}>=18'b001010000001011100) && ({row_reg, col_reg}<18'b001010000001100000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001010000001100000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001010000001100001) && ({row_reg, col_reg}<18'b001010000001100100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001010000001100100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001010000001100101) && ({row_reg, col_reg}<18'b001010000001101100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b001010000001101100) && ({row_reg, col_reg}<18'b001010000001101111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001010000001101111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001010000001110000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001010000001110001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001010000001110010)) color_data = 12'b011001010101;
		if(({row_reg, col_reg}>=18'b001010000001110011) && ({row_reg, col_reg}<18'b001010000001111001)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001010000001111001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b001010000001111010)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b001010000001111011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001010000001111100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001010000001111101) && ({row_reg, col_reg}<18'b001010000010000100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001010000010000100) && ({row_reg, col_reg}<18'b001010000010011100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b001010000010011100) && ({row_reg, col_reg}<18'b001010000010101100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001010000010101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001010000010101101)) color_data = 12'b011110001000;
		if(({row_reg, col_reg}==18'b001010000010101110)) color_data = 12'b011010001001;
		if(({row_reg, col_reg}==18'b001010000010101111)) color_data = 12'b100010011100;
		if(({row_reg, col_reg}==18'b001010000010110000)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}==18'b001010000010110001)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001010000010110010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001010000010110011) && ({row_reg, col_reg}<18'b001010000010110111)) color_data = 12'b011010101111;

		if(({row_reg, col_reg}>=18'b001010000010110111) && ({row_reg, col_reg}<18'b001010001001010011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001010001001010011) && ({row_reg, col_reg}<18'b001010001001010110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001010001001010110)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b001010001001010111) && ({row_reg, col_reg}<18'b001010001001011001)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b001010001001011001)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b001010001001011010)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b001010001001011011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001010001001011100) && ({row_reg, col_reg}<18'b001010001001100010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001010001001100010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001010001001100011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001010001001100100)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}>=18'b001010001001100101) && ({row_reg, col_reg}<18'b001010001001101100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001010001001101100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001010001001101101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001010001001101110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001010001001101111)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001010001001110000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001010001001110001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b001010001001110010) && ({row_reg, col_reg}<18'b001010001001110110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001010001001110110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001010001001110111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001010001001111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001010001001111001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b001010001001111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b001010001001111011) && ({row_reg, col_reg}<18'b001010001010000100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001010001010000100) && ({row_reg, col_reg}<18'b001010001010011100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001010001010011100)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b001010001010011101) && ({row_reg, col_reg}<18'b001010001010101100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001010001010101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001010001010101101)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==18'b001010001010101110)) color_data = 12'b011110001001;
		if(({row_reg, col_reg}==18'b001010001010101111)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b001010001010110000)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}==18'b001010001010110001)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001010001010110010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001010001010110011) && ({row_reg, col_reg}<18'b001010001010110110)) color_data = 12'b011010101111;

		if(({row_reg, col_reg}>=18'b001010001010110110) && ({row_reg, col_reg}<18'b001010010001010011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001010010001010011)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001010010001010100)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b001010010001010101) && ({row_reg, col_reg}<18'b001010010001010111)) color_data = 12'b011110011100;
		if(({row_reg, col_reg}==18'b001010010001010111)) color_data = 12'b100010011011;
		if(({row_reg, col_reg}==18'b001010010001011000)) color_data = 12'b100010011010;
		if(({row_reg, col_reg}==18'b001010010001011001)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b001010010001011010)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b001010010001011011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001010010001011100) && ({row_reg, col_reg}<18'b001010010001100000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b001010010001100000) && ({row_reg, col_reg}<18'b001010010001100010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001010010001100010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b001010010001100011) && ({row_reg, col_reg}<18'b001010010001100111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001010010001100111)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b001010010001101000) && ({row_reg, col_reg}<18'b001010010001101010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001010010001101010)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b001010010001101011) && ({row_reg, col_reg}<18'b001010010001101110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001010010001101110) && ({row_reg, col_reg}<18'b001010010001110000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b001010010001110000)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b001010010001110001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001010010001110010) && ({row_reg, col_reg}<18'b001010010001110110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001010010001110110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001010010001110111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001010010001111000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001010010001111001)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b001010010001111010)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b001010010001111011) && ({row_reg, col_reg}<18'b001010010001111110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001010010001111110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001010010001111111)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b001010010010000000) && ({row_reg, col_reg}<18'b001010010010000101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001010010010000101) && ({row_reg, col_reg}<18'b001010010010001100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001010010010001100)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b001010010010001101) && ({row_reg, col_reg}<18'b001010010010011001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001010010010011001)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001010010010011010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001010010010011011)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b001010010010011100) && ({row_reg, col_reg}<18'b001010010010101100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001010010010101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001010010010101101)) color_data = 12'b011110001000;
		if(({row_reg, col_reg}==18'b001010010010101110)) color_data = 12'b011110001001;
		if(({row_reg, col_reg}==18'b001010010010101111)) color_data = 12'b100010011011;
		if(({row_reg, col_reg}>=18'b001010010010110000) && ({row_reg, col_reg}<18'b001010010010110011)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001010010010110011)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}>=18'b001010010010110100) && ({row_reg, col_reg}<18'b001010010010110110)) color_data = 12'b011010101111;

		if(({row_reg, col_reg}>=18'b001010010010110110) && ({row_reg, col_reg}<18'b001010011001010010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001010011001010010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001010011001010011)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001010011001010100)) color_data = 12'b011110011100;
		if(({row_reg, col_reg}==18'b001010011001010101)) color_data = 12'b011010001010;
		if(({row_reg, col_reg}>=18'b001010011001010110) && ({row_reg, col_reg}<18'b001010011001011000)) color_data = 12'b011010001001;
		if(({row_reg, col_reg}==18'b001010011001011000)) color_data = 12'b011110001000;
		if(({row_reg, col_reg}==18'b001010011001011001)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}==18'b001010011001011010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001010011001011011) && ({row_reg, col_reg}<18'b001010011001100000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001010011001100000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==18'b001010011001100001)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001010011001100010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001010011001100011)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b001010011001100100) && ({row_reg, col_reg}<18'b001010011001100110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001010011001100110)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b001010011001100111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b001010011001101000) && ({row_reg, col_reg}<18'b001010011001101010)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b001010011001101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001010011001101011) && ({row_reg, col_reg}<18'b001010011001110100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001010011001110100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b001010011001110101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001010011001110110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b001010011001110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001010011001111000) && ({row_reg, col_reg}<18'b001010011010000100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001010011010000100)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b001010011010000101) && ({row_reg, col_reg}<18'b001010011010000111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001010011010000111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b001010011010001000) && ({row_reg, col_reg}<18'b001010011010011011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001010011010011011)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b001010011010011100) && ({row_reg, col_reg}<18'b001010011010100101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b001010011010100101) && ({row_reg, col_reg}<18'b001010011010101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001010011010101000) && ({row_reg, col_reg}<18'b001010011010101010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001010011010101010)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==18'b001010011010101011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001010011010101100)) color_data = 12'b011110000111;
		if(({row_reg, col_reg}==18'b001010011010101101)) color_data = 12'b011110001000;
		if(({row_reg, col_reg}==18'b001010011010101110)) color_data = 12'b011110001001;
		if(({row_reg, col_reg}==18'b001010011010101111)) color_data = 12'b100010011011;
		if(({row_reg, col_reg}==18'b001010011010110000)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b001010011010110001) && ({row_reg, col_reg}<18'b001010011010110011)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001010011010110011)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}==18'b001010011010110100)) color_data = 12'b011010101111;

		if(({row_reg, col_reg}>=18'b001010011010110101) && ({row_reg, col_reg}<18'b001010100001010001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001010100001010001)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001010100001010010) && ({row_reg, col_reg}<18'b001010100001010100)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001010100001010100)) color_data = 12'b011110011011;
		if(({row_reg, col_reg}==18'b001010100001010101)) color_data = 12'b011001111001;
		if(({row_reg, col_reg}>=18'b001010100001010110) && ({row_reg, col_reg}<18'b001010100001011000)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==18'b001010100001011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001010100001011001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b001010100001011010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001010100001011011) && ({row_reg, col_reg}<18'b001010100001100000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001010100001100000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001010100001100001)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001010100001100010)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001010100001100011) && ({row_reg, col_reg}<18'b001010100001100111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001010100001100111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b001010100001101000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001010100001101001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b001010100001101010) && ({row_reg, col_reg}<18'b001010100001110011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001010100001110011)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b001010100001110100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001010100001110101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b001010100001110110) && ({row_reg, col_reg}<18'b001010100001111100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001010100001111100)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b001010100001111101) && ({row_reg, col_reg}<18'b001010100001111111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001010100001111111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001010100010000000) && ({row_reg, col_reg}<18'b001010100010000100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001010100010000100)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b001010100010000101) && ({row_reg, col_reg}<18'b001010100010100101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001010100010100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001010100010100110) && ({row_reg, col_reg}<18'b001010100010101010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001010100010101010)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==18'b001010100010101011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001010100010101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001010100010101101)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==18'b001010100010101110)) color_data = 12'b011110001001;
		if(({row_reg, col_reg}==18'b001010100010101111)) color_data = 12'b100010011011;
		if(({row_reg, col_reg}>=18'b001010100010110000) && ({row_reg, col_reg}<18'b001010100010110010)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b001010100010110010) && ({row_reg, col_reg}<18'b001010100010110100)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001010100010110100)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}==18'b001010100010110101)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b001010100010110110) && ({row_reg, col_reg}<18'b001010101001001001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001010101001001001) && ({row_reg, col_reg}<18'b001010101001001100)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001010101001001100) && ({row_reg, col_reg}<18'b001010101001010000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001010101001010000) && ({row_reg, col_reg}<18'b001010101001010010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001010101001010010)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001010101001010011)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}==18'b001010101001010100)) color_data = 12'b011110011011;
		if(({row_reg, col_reg}==18'b001010101001010101)) color_data = 12'b011001111000;
		if(({row_reg, col_reg}==18'b001010101001010110)) color_data = 12'b011110001000;
		if(({row_reg, col_reg}==18'b001010101001010111)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b001010101001011000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001010101001011001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001010101001011010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001010101001011011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001010101001011100) && ({row_reg, col_reg}<18'b001010101001100000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001010101001100000)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==18'b001010101001100001)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001010101001100010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001010101001100011) && ({row_reg, col_reg}<18'b001010101001100111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001010101001100111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001010101001101000) && ({row_reg, col_reg}<18'b001010101001110101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001010101001110101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001010101001110110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001010101001110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001010101001111000) && ({row_reg, col_reg}<18'b001010101001111010)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b001010101001111010) && ({row_reg, col_reg}<18'b001010101010000100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001010101010000100)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b001010101010000101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001010101010000110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001010101010000111) && ({row_reg, col_reg}<18'b001010101010100101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001010101010100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001010101010100110) && ({row_reg, col_reg}<18'b001010101010101010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b001010101010101010) && ({row_reg, col_reg}<18'b001010101010101100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001010101010101100)) color_data = 12'b011110000111;
		if(({row_reg, col_reg}==18'b001010101010101101)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==18'b001010101010101110)) color_data = 12'b011110001001;
		if(({row_reg, col_reg}==18'b001010101010101111)) color_data = 12'b100010011011;
		if(({row_reg, col_reg}==18'b001010101010110000)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}==18'b001010101010110001)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b001010101010110010) && ({row_reg, col_reg}<18'b001010101010110110)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b001010101010110110) && ({row_reg, col_reg}<18'b001010110001001001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001010110001001001) && ({row_reg, col_reg}<18'b001010110001001101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001010110001001101) && ({row_reg, col_reg}<18'b001010110001010000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001010110001010000) && ({row_reg, col_reg}<18'b001010110001010010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001010110001010010)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001010110001010011)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}==18'b001010110001010100)) color_data = 12'b011110011011;
		if(({row_reg, col_reg}==18'b001010110001010101)) color_data = 12'b011001111000;
		if(({row_reg, col_reg}==18'b001010110001010110)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}>=18'b001010110001010111) && ({row_reg, col_reg}<18'b001010110001011001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001010110001011001)) color_data = 12'b101010011000;
		if(({row_reg, col_reg}==18'b001010110001011010)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==18'b001010110001011011)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b001010110001011100) && ({row_reg, col_reg}<18'b001010110001100010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001010110001100010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001010110001100011)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b001010110001100100) && ({row_reg, col_reg}<18'b001010110001100111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001010110001100111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001010110001101000) && ({row_reg, col_reg}<18'b001010110001110101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001010110001110101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b001010110001110110) && ({row_reg, col_reg}<18'b001010110001111010)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001010110001111010)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b001010110001111011) && ({row_reg, col_reg}<18'b001010110001111101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001010110001111101) && ({row_reg, col_reg}<18'b001010110001111111)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b001010110001111111) && ({row_reg, col_reg}<18'b001010110010000001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001010110010000001)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001010110010000010)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001010110010000011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b001010110010000100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b001010110010000101) && ({row_reg, col_reg}<18'b001010110010100101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b001010110010100101) && ({row_reg, col_reg}<18'b001010110010100111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001010110010100111) && ({row_reg, col_reg}<18'b001010110010101010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001010110010101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001010110010101011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001010110010101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001010110010101101)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==18'b001010110010101110)) color_data = 12'b011110001001;
		if(({row_reg, col_reg}==18'b001010110010101111)) color_data = 12'b100010011010;
		if(({row_reg, col_reg}>=18'b001010110010110000) && ({row_reg, col_reg}<18'b001010110010110010)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}>=18'b001010110010110010) && ({row_reg, col_reg}<18'b001010110010110100)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b001010110010110100) && ({row_reg, col_reg}<18'b001010110010110110)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b001010110010110110) && ({row_reg, col_reg}<18'b001010111001001001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001010111001001001) && ({row_reg, col_reg}<18'b001010111001001101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001010111001001101) && ({row_reg, col_reg}<18'b001010111001010010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001010111001010010)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001010111001010011)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}==18'b001010111001010100)) color_data = 12'b011110011011;
		if(({row_reg, col_reg}==18'b001010111001010101)) color_data = 12'b011001111000;
		if(({row_reg, col_reg}==18'b001010111001010110)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}>=18'b001010111001010111) && ({row_reg, col_reg}<18'b001010111001011001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001010111001011001)) color_data = 12'b101010011000;
		if(({row_reg, col_reg}==18'b001010111001011010)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}>=18'b001010111001011011) && ({row_reg, col_reg}<18'b001010111001011101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001010111001011101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001010111001011110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b001010111001011111)) color_data = 12'b100110001001;
		if(({row_reg, col_reg}==18'b001010111001100000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b001010111001100001) && ({row_reg, col_reg}<18'b001010111001100011)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b001010111001100011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001010111001100100) && ({row_reg, col_reg}<18'b001010111001100110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b001010111001100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001010111001100111) && ({row_reg, col_reg}<18'b001010111001110001)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b001010111001110001) && ({row_reg, col_reg}<18'b001010111001110011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001010111001110011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001010111001110100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001010111001110101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b001010111001110110) && ({row_reg, col_reg}<18'b001010111010000100)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b001010111010000100)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b001010111010000101) && ({row_reg, col_reg}<18'b001010111010000111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001010111010000111)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b001010111010001000) && ({row_reg, col_reg}<18'b001010111010101001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001010111010101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001010111010101010) && ({row_reg, col_reg}<18'b001010111010101100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b001010111010101100) && ({row_reg, col_reg}<18'b001010111010101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001010111010101110)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==18'b001010111010101111)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=18'b001010111010110000) && ({row_reg, col_reg}<18'b001010111010110010)) color_data = 12'b011110011010;
		if(({row_reg, col_reg}==18'b001010111010110010)) color_data = 12'b011110011011;
		if(({row_reg, col_reg}==18'b001010111010110011)) color_data = 12'b011010011100;
		if(({row_reg, col_reg}==18'b001010111010110100)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001010111010110101)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b001010111010110110) && ({row_reg, col_reg}<18'b001011000001001001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001011000001001001) && ({row_reg, col_reg}<18'b001011000001001101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001011000001001101) && ({row_reg, col_reg}<18'b001011000001010010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001011000001010010) && ({row_reg, col_reg}<18'b001011000001010100)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001011000001010100)) color_data = 12'b011110011011;
		if(({row_reg, col_reg}==18'b001011000001010101)) color_data = 12'b011001111000;
		if(({row_reg, col_reg}==18'b001011000001010110)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}>=18'b001011000001010111) && ({row_reg, col_reg}<18'b001011000001011001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001011000001011001)) color_data = 12'b101010011000;
		if(({row_reg, col_reg}>=18'b001011000001011010) && ({row_reg, col_reg}<18'b001011000001011101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001011000001011101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001011000001011110)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b001011000001011111) && ({row_reg, col_reg}<18'b001011000001100010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001011000001100010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001011000001100011) && ({row_reg, col_reg}<18'b001011000001110001)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b001011000001110001) && ({row_reg, col_reg}<18'b001011000001111101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001011000001111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001011000001111110) && ({row_reg, col_reg}<18'b001011000010101010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001011000010101010)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b001011000010101011) && ({row_reg, col_reg}<18'b001011000010101101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001011000010101101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b001011000010101110)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==18'b001011000010101111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001011000010110000)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==18'b001011000010110001)) color_data = 12'b011001111000;
		if(({row_reg, col_reg}==18'b001011000010110010)) color_data = 12'b011010001001;
		if(({row_reg, col_reg}==18'b001011000010110011)) color_data = 12'b011110011011;
		if(({row_reg, col_reg}==18'b001011000010110100)) color_data = 12'b011110011100;
		if(({row_reg, col_reg}==18'b001011000010110101)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b001011000010110110) && ({row_reg, col_reg}<18'b001011000010111000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001011000010111000)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b001011000010111001) && ({row_reg, col_reg}<18'b001011001001001000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001011001001001000) && ({row_reg, col_reg}<18'b001011001001001101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001011001001001101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001011001001001110) && ({row_reg, col_reg}<18'b001011001001010000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001011001001010000)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b001011001001010001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001011001001010010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001011001001010011)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001011001001010100)) color_data = 12'b011110011011;
		if(({row_reg, col_reg}==18'b001011001001010101)) color_data = 12'b011001111001;
		if(({row_reg, col_reg}==18'b001011001001010110)) color_data = 12'b011110001000;
		if(({row_reg, col_reg}==18'b001011001001010111)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}==18'b001011001001011000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001011001001011001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001011001001011010) && ({row_reg, col_reg}<18'b001011001001011101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001011001001011101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001011001001011110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b001011001001011111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001011001001100000) && ({row_reg, col_reg}<18'b001011001001100011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b001011001001100011) && ({row_reg, col_reg}<18'b001011001001110001)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b001011001001110001) && ({row_reg, col_reg}<18'b001011001010101010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b001011001010101010) && ({row_reg, col_reg}<18'b001011001010101111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001011001010101111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001011001010110000)) color_data = 12'b011110001000;
		if(({row_reg, col_reg}==18'b001011001010110001)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==18'b001011001010110010)) color_data = 12'b011001111001;
		if(({row_reg, col_reg}==18'b001011001010110011)) color_data = 12'b011110001010;
		if(({row_reg, col_reg}==18'b001011001010110100)) color_data = 12'b011110011100;
		if(({row_reg, col_reg}==18'b001011001010110101)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001011001010110110)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b001011001010110111) && ({row_reg, col_reg}<18'b001011010001001001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001011010001001001) && ({row_reg, col_reg}<18'b001011010001001100)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001011010001001100) && ({row_reg, col_reg}<18'b001011010001010010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001011010001010010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001011010001010011)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001011010001010100)) color_data = 12'b011110011011;
		if(({row_reg, col_reg}==18'b001011010001010101)) color_data = 12'b011001111001;
		if(({row_reg, col_reg}==18'b001011010001010110)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==18'b001011010001010111)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}==18'b001011010001011000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001011010001011001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001011010001011010) && ({row_reg, col_reg}<18'b001011010001011101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001011010001011101)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001011010001011110)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b001011010001011111) && ({row_reg, col_reg}<18'b001011010001100011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b001011010001100011) && ({row_reg, col_reg}<18'b001011010001110001)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b001011010001110001) && ({row_reg, col_reg}<18'b001011010010100100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001011010010100100)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b001011010010100101) && ({row_reg, col_reg}<18'b001011010010101010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001011010010101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001011010010101011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001011010010101100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b001011010010101101) && ({row_reg, col_reg}<18'b001011010010101111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b001011010010101111) && ({row_reg, col_reg}<18'b001011010010110001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001011010010110001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001011010010110010)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==18'b001011010010110011)) color_data = 12'b011110011010;
		if(({row_reg, col_reg}==18'b001011010010110100)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}==18'b001011010010110101)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}==18'b001011010010110110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001011010010110111) && ({row_reg, col_reg}<18'b001011010010111001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001011010010111001)) color_data = 12'b011010101111;

		if(({row_reg, col_reg}>=18'b001011010010111010) && ({row_reg, col_reg}<18'b001011011001001010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001011011001001010) && ({row_reg, col_reg}<18'b001011011001001101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001011011001001101) && ({row_reg, col_reg}<18'b001011011001010010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001011011001010010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001011011001010011)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001011011001010100)) color_data = 12'b011110011011;
		if(({row_reg, col_reg}==18'b001011011001010101)) color_data = 12'b011010001001;
		if(({row_reg, col_reg}>=18'b001011011001010110) && ({row_reg, col_reg}<18'b001011011001011000)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==18'b001011011001011000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b001011011001011001)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b001011011001011010)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==18'b001011011001011011)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001011011001011100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001011011001011101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001011011001011110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b001011011001011111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001011011001100000) && ({row_reg, col_reg}<18'b001011011001100010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001011011001100010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001011011001100011) && ({row_reg, col_reg}<18'b001011011001101101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001011011001101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001011011001101110) && ({row_reg, col_reg}<18'b001011011001110000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001011011001110000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001011011001110001) && ({row_reg, col_reg}<18'b001011011010100010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001011011010100010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001011011010100011)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b001011011010100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001011011010100101) && ({row_reg, col_reg}<18'b001011011010101010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001011011010101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001011011010101011) && ({row_reg, col_reg}<18'b001011011010101101)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b001011011010101101) && ({row_reg, col_reg}<18'b001011011010101111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001011011010101111)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==18'b001011011010110000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001011011010110001)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b001011011010110010)) color_data = 12'b011110001000;
		if(({row_reg, col_reg}==18'b001011011010110011)) color_data = 12'b100010011010;
		if(({row_reg, col_reg}==18'b001011011010110100)) color_data = 12'b011110011100;
		if(({row_reg, col_reg}==18'b001011011010110101)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001011011010110110)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b001011011010110111) && ({row_reg, col_reg}<18'b001011100001001000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001011100001001000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001011100001001001) && ({row_reg, col_reg}<18'b001011100001010000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001011100001010000) && ({row_reg, col_reg}<18'b001011100001010010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001011100001010010)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001011100001010011)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}==18'b001011100001010100)) color_data = 12'b011110011011;
		if(({row_reg, col_reg}==18'b001011100001010101)) color_data = 12'b011110001001;
		if(({row_reg, col_reg}==18'b001011100001010110)) color_data = 12'b011110001000;
		if(({row_reg, col_reg}==18'b001011100001010111)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==18'b001011100001011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001011100001011001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001011100001011010)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b001011100001011011)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b001011100001011100)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b001011100001011101)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b001011100001011110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b001011100001011111) && ({row_reg, col_reg}<18'b001011100001101100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001011100001101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001011100001101101) && ({row_reg, col_reg}<18'b001011100010100001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001011100010100001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001011100010100010) && ({row_reg, col_reg}<18'b001011100010100101)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b001011100010100101) && ({row_reg, col_reg}<18'b001011100010101011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001011100010101011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b001011100010101100) && ({row_reg, col_reg}<18'b001011100010101111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001011100010101111)) color_data = 12'b101010011000;
		if(({row_reg, col_reg}==18'b001011100010110000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001011100010110001) && ({row_reg, col_reg}<18'b001011100010110011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001011100010110011)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}==18'b001011100010110100)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b001011100010110101)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001011100010110110)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b001011100010110111) && ({row_reg, col_reg}<18'b001011101001010001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001011101001010001)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001011101001010010)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001011101001010011)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b001011101001010100)) color_data = 12'b011110011010;
		if(({row_reg, col_reg}==18'b001011101001010101)) color_data = 12'b011110001000;
		if(({row_reg, col_reg}==18'b001011101001010110)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==18'b001011101001010111)) color_data = 12'b011110000111;
		if(({row_reg, col_reg}>=18'b001011101001011000) && ({row_reg, col_reg}<18'b001011101001011100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001011101001011100) && ({row_reg, col_reg}<18'b001011101001011110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001011101001011110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001011101001011111)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}>=18'b001011101001100000) && ({row_reg, col_reg}<18'b001011101001101100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001011101001101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001011101001101101) && ({row_reg, col_reg}<18'b001011101010100001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b001011101010100001) && ({row_reg, col_reg}<18'b001011101010101011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001011101010101011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b001011101010101100) && ({row_reg, col_reg}<18'b001011101010101110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001011101010101110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b001011101010101111)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==18'b001011101010110000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001011101010110001)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==18'b001011101010110010)) color_data = 12'b101010111011;
		if(({row_reg, col_reg}==18'b001011101010110011)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b001011101010110100)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b001011101010110101)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001011101010110110)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b001011101010110111) && ({row_reg, col_reg}<18'b001011110001001110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001011110001001110)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b001011110001001111) && ({row_reg, col_reg}<18'b001011110001010001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001011110001010001) && ({row_reg, col_reg}<18'b001011110001010011)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001011110001010011)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b001011110001010100)) color_data = 12'b100010011010;
		if(({row_reg, col_reg}==18'b001011110001010101)) color_data = 12'b011110001000;
		if(({row_reg, col_reg}==18'b001011110001010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001011110001010111)) color_data = 12'b011110000111;
		if(({row_reg, col_reg}==18'b001011110001011000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b001011110001011001)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b001011110001011010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b001011110001011011) && ({row_reg, col_reg}<18'b001011110001011110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001011110001011110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b001011110001011111) && ({row_reg, col_reg}<18'b001011110001101100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001011110001101100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b001011110001101101) && ({row_reg, col_reg}<18'b001011110010100001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b001011110010100001) && ({row_reg, col_reg}<18'b001011110010101011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001011110010101011)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b001011110010101100) && ({row_reg, col_reg}<18'b001011110010101111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001011110010101111)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==18'b001011110010110000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001011110010110001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001011110010110010)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b001011110010110011)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b001011110010110100)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b001011110010110101)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001011110010110110)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b001011110010110111) && ({row_reg, col_reg}<18'b001011111001001000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001011111001001000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001011111001001001) && ({row_reg, col_reg}<18'b001011111001001110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001011111001001110) && ({row_reg, col_reg}<18'b001011111001010000)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b001011111001010000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001011111001010001)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001011111001010010)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}==18'b001011111001010011)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==18'b001011111001010100)) color_data = 12'b100010011010;
		if(({row_reg, col_reg}==18'b001011111001010101)) color_data = 12'b011110001000;
		if(({row_reg, col_reg}==18'b001011111001010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001011111001010111) && ({row_reg, col_reg}<18'b001011111001011010)) color_data = 12'b011110000111;
		if(({row_reg, col_reg}==18'b001011111001011010)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b001011111001011011) && ({row_reg, col_reg}<18'b001011111001011101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001011111001011101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001011111001011110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b001011111001011111) && ({row_reg, col_reg}<18'b001011111001101100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001011111001101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001011111001101101) && ({row_reg, col_reg}<18'b001011111010100001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b001011111010100001) && ({row_reg, col_reg}<18'b001011111010101011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001011111010101011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001011111010101100) && ({row_reg, col_reg}<18'b001011111010101111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001011111010101111)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}>=18'b001011111010110000) && ({row_reg, col_reg}<18'b001011111010110010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001011111010110010)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b001011111010110011)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b001011111010110100)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}>=18'b001011111010110101) && ({row_reg, col_reg}<18'b001011111010110111)) color_data = 12'b011110101101;

		if(({row_reg, col_reg}>=18'b001011111010110111) && ({row_reg, col_reg}<18'b001100000001000010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001100000001000010) && ({row_reg, col_reg}<18'b001100000001000101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001100000001000101) && ({row_reg, col_reg}<18'b001100000001001000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001100000001001000) && ({row_reg, col_reg}<18'b001100000001001011)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b001100000001001011) && ({row_reg, col_reg}<18'b001100000001001101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001100000001001101) && ({row_reg, col_reg}<18'b001100000001010000)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b001100000001010000) && ({row_reg, col_reg}<18'b001100000001010010)) color_data = 12'b011110011010;
		if(({row_reg, col_reg}==18'b001100000001010010)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}==18'b001100000001010011)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}==18'b001100000001010100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b001100000001010101) && ({row_reg, col_reg}<18'b001100000001011001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b001100000001011001) && ({row_reg, col_reg}<18'b001100000001011101)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b001100000001011101) && ({row_reg, col_reg}<18'b001100000001101100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001100000001101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001100000001101101) && ({row_reg, col_reg}<18'b001100000010010111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001100000010010111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001100000010011000)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b001100000010011001) && ({row_reg, col_reg}<18'b001100000010100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001100000010100000) && ({row_reg, col_reg}<18'b001100000010101110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001100000010101110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b001100000010101111)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b001100000010110000) && ({row_reg, col_reg}<18'b001100000010110010)) color_data = 12'b101010111010;
		if(({row_reg, col_reg}==18'b001100000010110010)) color_data = 12'b100110111011;
		if(({row_reg, col_reg}==18'b001100000010110011)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b001100000010110100)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001100000010110101)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}>=18'b001100000010110110) && ({row_reg, col_reg}<18'b001100000010111010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001100000010111010) && ({row_reg, col_reg}<18'b001100000010111110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001100000010111110) && ({row_reg, col_reg}<18'b001100000011010100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001100000011010100) && ({row_reg, col_reg}<18'b001100000011010110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001100000011010110) && ({row_reg, col_reg}<18'b001100000011101111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001100000011101111)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b001100000011110000) && ({row_reg, col_reg}<18'b001100001001000010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001100001001000010) && ({row_reg, col_reg}<18'b001100001001000101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001100001001000101) && ({row_reg, col_reg}<18'b001100001001001000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001100001001001000) && ({row_reg, col_reg}<18'b001100001001001011)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b001100001001001011) && ({row_reg, col_reg}<18'b001100001001001101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001100001001001101)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}==18'b001100001001001110)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001100001001001111)) color_data = 12'b011010011100;
		if(({row_reg, col_reg}==18'b001100001001010000)) color_data = 12'b011010001001;
		if(({row_reg, col_reg}==18'b001100001001010001)) color_data = 12'b011010001000;
		if(({row_reg, col_reg}==18'b001100001001010010)) color_data = 12'b011001111000;
		if(({row_reg, col_reg}==18'b001100001001010011)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}>=18'b001100001001010100) && ({row_reg, col_reg}<18'b001100001001010111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001100001001010111)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b001100001001011000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001100001001011001)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b001100001001011010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001100001001011011)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b001100001001011100) && ({row_reg, col_reg}<18'b001100001001101100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001100001001101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001100001001101101) && ({row_reg, col_reg}<18'b001100001010010111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001100001010010111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b001100001010011000) && ({row_reg, col_reg}<18'b001100001010101110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001100001010101110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b001100001010101111) && ({row_reg, col_reg}<18'b001100001010110001)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001100001010110001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001100001010110010)) color_data = 12'b100110111011;
		if(({row_reg, col_reg}==18'b001100001010110011)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}>=18'b001100001010110100) && ({row_reg, col_reg}<18'b001100001010110110)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b001100001010110110) && ({row_reg, col_reg}<18'b001100001010111010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001100001010111010) && ({row_reg, col_reg}<18'b001100001010111101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001100001010111101) && ({row_reg, col_reg}<18'b001100001011011111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001100001011011111)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001100001011100000) && ({row_reg, col_reg}<18'b001100001011101111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001100001011101111)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b001100001011110000) && ({row_reg, col_reg}<18'b001100010001000011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001100010001000011) && ({row_reg, col_reg}<18'b001100010001000101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001100010001000101) && ({row_reg, col_reg}<18'b001100010001001001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001100010001001001)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b001100010001001010) && ({row_reg, col_reg}<18'b001100010001001101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001100010001001101) && ({row_reg, col_reg}<18'b001100010001001111)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001100010001001111)) color_data = 12'b011110011100;
		if(({row_reg, col_reg}>=18'b001100010001010000) && ({row_reg, col_reg}<18'b001100010001010010)) color_data = 12'b011010001001;
		if(({row_reg, col_reg}==18'b001100010001010010)) color_data = 12'b011110001000;
		if(({row_reg, col_reg}==18'b001100010001010011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001100010001010100) && ({row_reg, col_reg}<18'b001100010001011001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001100010001011001)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b001100010001011010) && ({row_reg, col_reg}<18'b001100010001101100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001100010001101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001100010001101101) && ({row_reg, col_reg}<18'b001100010010010111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001100010010010111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b001100010010011000) && ({row_reg, col_reg}<18'b001100010010101110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001100010010101110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b001100010010101111) && ({row_reg, col_reg}<18'b001100010010110001)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001100010010110001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001100010010110010)) color_data = 12'b100110111011;
		if(({row_reg, col_reg}==18'b001100010010110011)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}>=18'b001100010010110100) && ({row_reg, col_reg}<18'b001100010010110110)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001100010010110110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001100010010110111) && ({row_reg, col_reg}<18'b001100010010111011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001100010010111011)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001100010010111100) && ({row_reg, col_reg}<18'b001100010011001000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001100010011001000)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b001100010011001001) && ({row_reg, col_reg}<18'b001100010011011110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001100010011011110) && ({row_reg, col_reg}<18'b001100010011100000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001100010011100000) && ({row_reg, col_reg}<18'b001100010011100011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001100010011100011) && ({row_reg, col_reg}<18'b001100010011100110)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b001100010011100110) && ({row_reg, col_reg}<18'b001100011001001101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001100011001001101) && ({row_reg, col_reg}<18'b001100011001001111)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001100011001001111)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}==18'b001100011001010000)) color_data = 12'b011010001000;
		if(({row_reg, col_reg}>=18'b001100011001010001) && ({row_reg, col_reg}<18'b001100011001010011)) color_data = 12'b011110001000;
		if(({row_reg, col_reg}==18'b001100011001010011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b001100011001010100) && ({row_reg, col_reg}<18'b001100011001010111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001100011001010111)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b001100011001011000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001100011001011001)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b001100011001011010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b001100011001011011) && ({row_reg, col_reg}<18'b001100011001101100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001100011001101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001100011001101101) && ({row_reg, col_reg}<18'b001100011010010111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001100011010010111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b001100011010011000) && ({row_reg, col_reg}<18'b001100011010101110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001100011010101110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b001100011010101111)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b001100011010110000) && ({row_reg, col_reg}<18'b001100011010110010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001100011010110010)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b001100011010110011)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==18'b001100011010110100)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}==18'b001100011010110101)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b001100011010110110) && ({row_reg, col_reg}<18'b001100011011000000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001100011011000000) && ({row_reg, col_reg}<18'b001100011011000100)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001100011011000100) && ({row_reg, col_reg}<18'b001100011011000110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001100011011000110) && ({row_reg, col_reg}<18'b001100011011001100)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b001100011011001100) && ({row_reg, col_reg}<18'b001100011011011101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001100011011011101) && ({row_reg, col_reg}<18'b001100011011100000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001100011011100000) && ({row_reg, col_reg}<18'b001100011011100010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001100011011100010) && ({row_reg, col_reg}<18'b001100011011100111)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b001100011011100111) && ({row_reg, col_reg}<18'b001100100001001101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001100100001001101) && ({row_reg, col_reg}<18'b001100100001001111)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001100100001001111)) color_data = 12'b011110011100;
		if(({row_reg, col_reg}==18'b001100100001010000)) color_data = 12'b011010001000;
		if(({row_reg, col_reg}==18'b001100100001010001)) color_data = 12'b011110001000;
		if(({row_reg, col_reg}==18'b001100100001010010)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}>=18'b001100100001010011) && ({row_reg, col_reg}<18'b001100100001010101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001100100001010101)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}>=18'b001100100001010110) && ({row_reg, col_reg}<18'b001100100001011001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001100100001011001)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b001100100001011010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b001100100001011011) && ({row_reg, col_reg}<18'b001100100001101100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001100100001101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001100100001101101) && ({row_reg, col_reg}<18'b001100100010010011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001100100010010011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001100100010010100) && ({row_reg, col_reg}<18'b001100100010010111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001100100010010111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b001100100010011000) && ({row_reg, col_reg}<18'b001100100010101110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001100100010101110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b001100100010101111)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001100100010110000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001100100010110001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001100100010110010)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b001100100010110011)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==18'b001100100010110100)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}==18'b001100100010110101)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001100100010110110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001100100010110111) && ({row_reg, col_reg}<18'b001100100011000000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001100100011000000) && ({row_reg, col_reg}<18'b001100100011000101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001100100011000101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001100100011000110) && ({row_reg, col_reg}<18'b001100100011001110)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b001100100011001110) && ({row_reg, col_reg}<18'b001100100011010110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001100100011010110) && ({row_reg, col_reg}<18'b001100100011011000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001100100011011000) && ({row_reg, col_reg}<18'b001100100011011101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001100100011011101) && ({row_reg, col_reg}<18'b001100100011100000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001100100011100000) && ({row_reg, col_reg}<18'b001100100011100010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001100100011100010) && ({row_reg, col_reg}<18'b001100100011101000)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b001100100011101000) && ({row_reg, col_reg}<18'b001100101001000111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001100101001000111) && ({row_reg, col_reg}<18'b001100101001001001)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001100101001001001) && ({row_reg, col_reg}<18'b001100101001001101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001100101001001101) && ({row_reg, col_reg}<18'b001100101001001111)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001100101001001111)) color_data = 12'b011110011011;
		if(({row_reg, col_reg}>=18'b001100101001010000) && ({row_reg, col_reg}<18'b001100101001010010)) color_data = 12'b011110001000;
		if(({row_reg, col_reg}==18'b001100101001010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001100101001010011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001100101001010100)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}>=18'b001100101001010101) && ({row_reg, col_reg}<18'b001100101001010111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b001100101001010111) && ({row_reg, col_reg}<18'b001100101001011001)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b001100101001011001)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001100101001011010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b001100101001011011) && ({row_reg, col_reg}<18'b001100101001101100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001100101001101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001100101001101101) && ({row_reg, col_reg}<18'b001100101010010010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001100101010010010)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b001100101010010011) && ({row_reg, col_reg}<18'b001100101010010101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b001100101010010101) && ({row_reg, col_reg}<18'b001100101010010111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b001100101010010111) && ({row_reg, col_reg}<18'b001100101010101110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001100101010101110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b001100101010101111)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001100101010110000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001100101010110001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001100101010110010)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b001100101010110011)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==18'b001100101010110100)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}==18'b001100101010110101)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001100101010110110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001100101010110111) && ({row_reg, col_reg}<18'b001100101011000000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001100101011000000) && ({row_reg, col_reg}<18'b001100101011000110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001100101011000110) && ({row_reg, col_reg}<18'b001100101011001001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001100101011001001) && ({row_reg, col_reg}<18'b001100101011010000)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b001100101011010000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001100101011010001) && ({row_reg, col_reg}<18'b001100101011010101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001100101011010101) && ({row_reg, col_reg}<18'b001100101011011010)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}==18'b001100101011011010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001100101011011011)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001100101011011100) && ({row_reg, col_reg}<18'b001100101011011110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001100101011011110) && ({row_reg, col_reg}<18'b001100101011100000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001100101011100000) && ({row_reg, col_reg}<18'b001100101011100010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001100101011100010) && ({row_reg, col_reg}<18'b001100101011101001)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b001100101011101001) && ({row_reg, col_reg}<18'b001100110001000111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001100110001000111) && ({row_reg, col_reg}<18'b001100110001001001)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001100110001001001) && ({row_reg, col_reg}<18'b001100110001001101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001100110001001101) && ({row_reg, col_reg}<18'b001100110001001111)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001100110001001111)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}>=18'b001100110001010000) && ({row_reg, col_reg}<18'b001100110001010010)) color_data = 12'b011110001000;
		if(({row_reg, col_reg}==18'b001100110001010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001100110001010011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001100110001010100)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}>=18'b001100110001010101) && ({row_reg, col_reg}<18'b001100110001011010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001100110001011010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b001100110001011011) && ({row_reg, col_reg}<18'b001100110001101100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001100110001101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001100110001101101) && ({row_reg, col_reg}<18'b001100110010010010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001100110010010010)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b001100110010010011) && ({row_reg, col_reg}<18'b001100110010101110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001100110010101110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b001100110010101111)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001100110010110000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001100110010110001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001100110010110010)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b001100110010110011)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==18'b001100110010110100)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}==18'b001100110010110101)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001100110010110110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001100110010110111) && ({row_reg, col_reg}<18'b001100110011000000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001100110011000000) && ({row_reg, col_reg}<18'b001100110011010101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001100110011010101) && ({row_reg, col_reg}<18'b001100110011011011)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}>=18'b001100110011011011) && ({row_reg, col_reg}<18'b001100110011100011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001100110011100011) && ({row_reg, col_reg}<18'b001100110011101001)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b001100110011101001) && ({row_reg, col_reg}<18'b001100111001000000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001100111001000000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001100111001000001) && ({row_reg, col_reg}<18'b001100111001000110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001100111001000110) && ({row_reg, col_reg}<18'b001100111001001000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001100111001001000) && ({row_reg, col_reg}<18'b001100111001001101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001100111001001101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001100111001001110)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001100111001001111)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}>=18'b001100111001010000) && ({row_reg, col_reg}<18'b001100111001010011)) color_data = 12'b011110001000;
		if(({row_reg, col_reg}>=18'b001100111001010011) && ({row_reg, col_reg}<18'b001100111001010101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b001100111001010101) && ({row_reg, col_reg}<18'b001100111001101100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001100111001101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001100111001101101) && ({row_reg, col_reg}<18'b001100111010010010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001100111010010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001100111010010011) && ({row_reg, col_reg}<18'b001100111010101110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001100111010101110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b001100111010101111)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001100111010110000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001100111010110001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001100111010110010)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b001100111010110011)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==18'b001100111010110100)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}==18'b001100111010110101)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001100111010110110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001100111010110111) && ({row_reg, col_reg}<18'b001100111011000000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001100111011000000)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b001100111011000001) && ({row_reg, col_reg}<18'b001100111011000011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001100111011000011) && ({row_reg, col_reg}<18'b001100111011000111)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001100111011000111) && ({row_reg, col_reg}<18'b001100111011001100)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b001100111011001100) && ({row_reg, col_reg}<18'b001100111011010000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001100111011010000) && ({row_reg, col_reg}<18'b001100111011010010)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b001100111011010010) && ({row_reg, col_reg}<18'b001100111011011001)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001100111011011001)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}==18'b001100111011011010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001100111011011011) && ({row_reg, col_reg}<18'b001100111011100110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001100111011100110) && ({row_reg, col_reg}<18'b001100111011101010)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b001100111011101010) && ({row_reg, col_reg}<18'b001101000001000000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001101000001000000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001101000001000001) && ({row_reg, col_reg}<18'b001101000001000110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001101000001000110) && ({row_reg, col_reg}<18'b001101000001001000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001101000001001000) && ({row_reg, col_reg}<18'b001101000001001011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001101000001001011)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b001101000001001100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001101000001001101) && ({row_reg, col_reg}<18'b001101000001001111)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001101000001001111)) color_data = 12'b011110011100;
		if(({row_reg, col_reg}==18'b001101000001010000)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==18'b001101000001010001)) color_data = 12'b011110001000;
		if(({row_reg, col_reg}==18'b001101000001010010)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==18'b001101000001010011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001101000001010100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b001101000001010101) && ({row_reg, col_reg}<18'b001101000001101100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001101000001101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001101000001101101) && ({row_reg, col_reg}<18'b001101000010010010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001101000010010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001101000010010011) && ({row_reg, col_reg}<18'b001101000010101110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001101000010101110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b001101000010101111)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001101000010110000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001101000010110001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001101000010110010)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b001101000010110011)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==18'b001101000010110100)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}==18'b001101000010110101)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b001101000010110110) && ({row_reg, col_reg}<18'b001101000010111000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001101000010111000) && ({row_reg, col_reg}<18'b001101000010111011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001101000010111011)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001101000010111100) && ({row_reg, col_reg}<18'b001101000011000000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001101000011000000) && ({row_reg, col_reg}<18'b001101000011000010)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b001101000011000010) && ({row_reg, col_reg}<18'b001101000011000100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001101000011000100)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001101000011000101) && ({row_reg, col_reg}<18'b001101000011001000)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b001101000011001000) && ({row_reg, col_reg}<18'b001101000011001010)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}>=18'b001101000011001010) && ({row_reg, col_reg}<18'b001101000011001100)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}>=18'b001101000011001100) && ({row_reg, col_reg}<18'b001101000011010000)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}==18'b001101000011010000)) color_data = 12'b100010011100;
		if(({row_reg, col_reg}>=18'b001101000011010001) && ({row_reg, col_reg}<18'b001101000011010101)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}>=18'b001101000011010101) && ({row_reg, col_reg}<18'b001101000011011000)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b001101000011011000) && ({row_reg, col_reg}<18'b001101000011011100)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001101000011011100) && ({row_reg, col_reg}<18'b001101000011011111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001101000011011111)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b001101000011100000) && ({row_reg, col_reg}<18'b001101000011101000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001101000011101000) && ({row_reg, col_reg}<18'b001101000011101011)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b001101000011101011) && ({row_reg, col_reg}<18'b001101001001000000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001101001001000000) && ({row_reg, col_reg}<18'b001101001001000010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001101001001000010) && ({row_reg, col_reg}<18'b001101001001000110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001101001001000110) && ({row_reg, col_reg}<18'b001101001001001000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001101001001001000) && ({row_reg, col_reg}<18'b001101001001001010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001101001001001010) && ({row_reg, col_reg}<18'b001101001001001100)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b001101001001001100)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}>=18'b001101001001001101) && ({row_reg, col_reg}<18'b001101001001001111)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001101001001001111)) color_data = 12'b011110011011;
		if(({row_reg, col_reg}==18'b001101001001010000)) color_data = 12'b011001111000;
		if(({row_reg, col_reg}==18'b001101001001010001)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}>=18'b001101001001010010) && ({row_reg, col_reg}<18'b001101001001010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001101001001010100) && ({row_reg, col_reg}<18'b001101001001101100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001101001001101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001101001001101101) && ({row_reg, col_reg}<18'b001101001010001110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001101001010001110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001101001010001111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b001101001010010000) && ({row_reg, col_reg}<18'b001101001010010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001101001010010010) && ({row_reg, col_reg}<18'b001101001010101110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001101001010101110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b001101001010101111)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b001101001010110000) && ({row_reg, col_reg}<18'b001101001010110010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001101001010110010)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b001101001010110011)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==18'b001101001010110100)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}==18'b001101001010110101)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b001101001010110110) && ({row_reg, col_reg}<18'b001101001010111000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001101001010111000) && ({row_reg, col_reg}<18'b001101001010111011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001101001010111011)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001101001010111100) && ({row_reg, col_reg}<18'b001101001010111110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001101001010111110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001101001010111111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001101001011000000) && ({row_reg, col_reg}<18'b001101001011000010)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b001101001011000010) && ({row_reg, col_reg}<18'b001101001011000100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001101001011000100)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001101001011000101) && ({row_reg, col_reg}<18'b001101001011000111)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001101001011000111)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}>=18'b001101001011001000) && ({row_reg, col_reg}<18'b001101001011001011)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}>=18'b001101001011001011) && ({row_reg, col_reg}<18'b001101001011010101)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}>=18'b001101001011010101) && ({row_reg, col_reg}<18'b001101001011011000)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b001101001011011000)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}>=18'b001101001011011001) && ({row_reg, col_reg}<18'b001101001011011100)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b001101001011011100) && ({row_reg, col_reg}<18'b001101001011011110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001101001011011110) && ({row_reg, col_reg}<18'b001101001011100000)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b001101001011100000) && ({row_reg, col_reg}<18'b001101001011101001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001101001011101001) && ({row_reg, col_reg}<18'b001101001011101100)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b001101001011101100) && ({row_reg, col_reg}<18'b001101010001000000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001101010001000000) && ({row_reg, col_reg}<18'b001101010001000010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001101010001000010) && ({row_reg, col_reg}<18'b001101010001000110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001101010001000110) && ({row_reg, col_reg}<18'b001101010001001000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001101010001001000) && ({row_reg, col_reg}<18'b001101010001001100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001101010001001100)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001101010001001101)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001101010001001110)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}==18'b001101010001001111)) color_data = 12'b011110011011;
		if(({row_reg, col_reg}>=18'b001101010001010000) && ({row_reg, col_reg}<18'b001101010001010010)) color_data = 12'b011001111000;
		if(({row_reg, col_reg}==18'b001101010001010010)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}>=18'b001101010001010011) && ({row_reg, col_reg}<18'b001101010001101100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001101010001101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001101010001101101) && ({row_reg, col_reg}<18'b001101010010001101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001101010010001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001101010010001110) && ({row_reg, col_reg}<18'b001101010010101110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001101010010101110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b001101010010101111)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b001101010010110000) && ({row_reg, col_reg}<18'b001101010010110010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001101010010110010)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b001101010010110011)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==18'b001101010010110100)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}==18'b001101010010110101)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b001101010010110110) && ({row_reg, col_reg}<18'b001101010010111000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001101010010111000) && ({row_reg, col_reg}<18'b001101010010111011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001101010010111011) && ({row_reg, col_reg}<18'b001101010011000000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001101010011000000) && ({row_reg, col_reg}<18'b001101010011000010)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b001101010011000010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001101010011000011)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001101010011000100) && ({row_reg, col_reg}<18'b001101010011000110)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001101010011000110)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}==18'b001101010011000111)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}>=18'b001101010011001000) && ({row_reg, col_reg}<18'b001101010011001010)) color_data = 12'b100110111100;
		if(({row_reg, col_reg}==18'b001101010011001010)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}>=18'b001101010011001011) && ({row_reg, col_reg}<18'b001101010011010100)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}>=18'b001101010011010100) && ({row_reg, col_reg}<18'b001101010011010110)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}>=18'b001101010011010110) && ({row_reg, col_reg}<18'b001101010011011001)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}==18'b001101010011011001)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b001101010011011010)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}>=18'b001101010011011011) && ({row_reg, col_reg}<18'b001101010011011101)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b001101010011011101) && ({row_reg, col_reg}<18'b001101010011011111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001101010011011111)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b001101010011100000) && ({row_reg, col_reg}<18'b001101010011101010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001101010011101010) && ({row_reg, col_reg}<18'b001101010011101100)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b001101010011101100) && ({row_reg, col_reg}<18'b001101011001000000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001101011001000000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001101011001000001) && ({row_reg, col_reg}<18'b001101011001000110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001101011001000110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001101011001000111) && ({row_reg, col_reg}<18'b001101011001001011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001101011001001011)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001101011001001100)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001101011001001101)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}==18'b001101011001001110)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b001101011001001111)) color_data = 12'b011110011011;
		if(({row_reg, col_reg}==18'b001101011001010000)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}>=18'b001101011001010001) && ({row_reg, col_reg}<18'b001101011001010011)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}==18'b001101011001010011)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b001101011001010100) && ({row_reg, col_reg}<18'b001101011001101100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001101011001101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001101011001101101) && ({row_reg, col_reg}<18'b001101011010001101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001101011010001101)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b001101011010001110) && ({row_reg, col_reg}<18'b001101011010101110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001101011010101110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b001101011010101111)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001101011010110000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001101011010110001) && ({row_reg, col_reg}<18'b001101011010110011)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b001101011010110011)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==18'b001101011010110100)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b001101011010110101)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b001101011010110110) && ({row_reg, col_reg}<18'b001101011010111000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001101011010111000) && ({row_reg, col_reg}<18'b001101011010111010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001101011010111010) && ({row_reg, col_reg}<18'b001101011010111100)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001101011010111100) && ({row_reg, col_reg}<18'b001101011010111110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001101011010111110) && ({row_reg, col_reg}<18'b001101011011000000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001101011011000000)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b001101011011000001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001101011011000010) && ({row_reg, col_reg}<18'b001101011011000100)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001101011011000100) && ({row_reg, col_reg}<18'b001101011011000110)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001101011011000110)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b001101011011000111)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==18'b001101011011001000)) color_data = 12'b101010111100;
		if(({row_reg, col_reg}==18'b001101011011001001)) color_data = 12'b101010111011;
		if(({row_reg, col_reg}>=18'b001101011011001010) && ({row_reg, col_reg}<18'b001101011011001100)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}>=18'b001101011011001100) && ({row_reg, col_reg}<18'b001101011011010000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001101011011010000)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}>=18'b001101011011010001) && ({row_reg, col_reg}<18'b001101011011010110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001101011011010110) && ({row_reg, col_reg}<18'b001101011011011000)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==18'b001101011011011000)) color_data = 12'b100010101010;
		if(({row_reg, col_reg}>=18'b001101011011011001) && ({row_reg, col_reg}<18'b001101011011011011)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}==18'b001101011011011011)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}>=18'b001101011011011100) && ({row_reg, col_reg}<18'b001101011011011110)) color_data = 12'b011110101101;

		if(({row_reg, col_reg}>=18'b001101011011011110) && ({row_reg, col_reg}<18'b001101100001000000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001101100001000000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001101100001000001) && ({row_reg, col_reg}<18'b001101100001000110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001101100001000110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001101100001000111) && ({row_reg, col_reg}<18'b001101100001001011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001101100001001011) && ({row_reg, col_reg}<18'b001101100001001101)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001101100001001101)) color_data = 12'b100010011100;
		if(({row_reg, col_reg}==18'b001101100001001110)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==18'b001101100001001111)) color_data = 12'b100010011010;
		if(({row_reg, col_reg}>=18'b001101100001010000) && ({row_reg, col_reg}<18'b001101100001010011)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}>=18'b001101100001010011) && ({row_reg, col_reg}<18'b001101100001101100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001101100001101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001101100001101101) && ({row_reg, col_reg}<18'b001101100010001110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001101100010001110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b001101100010001111) && ({row_reg, col_reg}<18'b001101100010101110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001101100010101110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b001101100010101111)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001101100010110000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001101100010110001) && ({row_reg, col_reg}<18'b001101100010110011)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b001101100010110011)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==18'b001101100010110100)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b001101100010110101)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b001101100010110110) && ({row_reg, col_reg}<18'b001101100010111000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001101100010111000) && ({row_reg, col_reg}<18'b001101100010111010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001101100010111010) && ({row_reg, col_reg}<18'b001101100010111100)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001101100010111100) && ({row_reg, col_reg}<18'b001101100010111110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001101100010111110) && ({row_reg, col_reg}<18'b001101100011000000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001101100011000000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001101100011000001) && ({row_reg, col_reg}<18'b001101100011000011)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001101100011000011)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001101100011000100)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}==18'b001101100011000101)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b001101100011000110)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==18'b001101100011000111)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}>=18'b001101100011001000) && ({row_reg, col_reg}<18'b001101100011001010)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}>=18'b001101100011001010) && ({row_reg, col_reg}<18'b001101100011001101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001101100011001101) && ({row_reg, col_reg}<18'b001101100011010011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b001101100011010011) && ({row_reg, col_reg}<18'b001101100011010110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001101100011010110)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001101100011010111)) color_data = 12'b100110101001;
		if(({row_reg, col_reg}>=18'b001101100011011000) && ({row_reg, col_reg}<18'b001101100011011010)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}>=18'b001101100011011010) && ({row_reg, col_reg}<18'b001101100011011100)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}==18'b001101100011011100)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}>=18'b001101100011011101) && ({row_reg, col_reg}<18'b001101100011011111)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b001101100011011111) && ({row_reg, col_reg}<18'b001101100011100001)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b001101100011100001) && ({row_reg, col_reg}<18'b001101101001000000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001101101001000000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001101101001000001) && ({row_reg, col_reg}<18'b001101101001000110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001101101001000110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001101101001000111) && ({row_reg, col_reg}<18'b001101101001001010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001101101001001010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001101101001001011)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001101101001001100)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b001101101001001101)) color_data = 12'b100010011011;
		if(({row_reg, col_reg}==18'b001101101001001110)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b001101101001001111)) color_data = 12'b100010011010;
		if(({row_reg, col_reg}==18'b001101101001010000)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}>=18'b001101101001010001) && ({row_reg, col_reg}<18'b001101101001010011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b001101101001010011) && ({row_reg, col_reg}<18'b001101101001101100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001101101001101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001101101001101101) && ({row_reg, col_reg}<18'b001101101010001101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001101101010001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001101101010001110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b001101101010001111) && ({row_reg, col_reg}<18'b001101101010101110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001101101010101110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b001101101010101111)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001101101010110000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001101101010110001) && ({row_reg, col_reg}<18'b001101101010110011)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b001101101010110011)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==18'b001101101010110100)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b001101101010110101)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b001101101010110110) && ({row_reg, col_reg}<18'b001101101010111000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001101101010111000) && ({row_reg, col_reg}<18'b001101101010111110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001101101010111110) && ({row_reg, col_reg}<18'b001101101011000001)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001101101011000001) && ({row_reg, col_reg}<18'b001101101011000011)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001101101011000011)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}==18'b001101101011000100)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b001101101011000101)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}==18'b001101101011000110)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}>=18'b001101101011000111) && ({row_reg, col_reg}<18'b001101101011001001)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}>=18'b001101101011001001) && ({row_reg, col_reg}<18'b001101101011010100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b001101101011010100) && ({row_reg, col_reg}<18'b001101101011010110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001101101011010110)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001101101011010111)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}>=18'b001101101011011000) && ({row_reg, col_reg}<18'b001101101011011010)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==18'b001101101011011010)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b001101101011011011)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}==18'b001101101011011100)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b001101101011011101)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}>=18'b001101101011011110) && ({row_reg, col_reg}<18'b001101101011100000)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b001101101011100000) && ({row_reg, col_reg}<18'b001101101011100011)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b001101101011100011) && ({row_reg, col_reg}<18'b001101110001000110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001101110001000110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001101110001000111) && ({row_reg, col_reg}<18'b001101110001001010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001101110001001010)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001101110001001011)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}==18'b001101110001001100)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==18'b001101110001001101)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b001101110001001110)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b001101110001001111)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}==18'b001101110001010000)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==18'b001101110001010001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b001101110001010010) && ({row_reg, col_reg}<18'b001101110001101100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001101110001101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001101110001101101) && ({row_reg, col_reg}<18'b001101110010001001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001101110010001001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001101110010001010) && ({row_reg, col_reg}<18'b001101110010101110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001101110010101110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b001101110010101111)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001101110010110000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001101110010110001) && ({row_reg, col_reg}<18'b001101110010110011)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b001101110010110011)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==18'b001101110010110100)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b001101110010110101)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b001101110010110110) && ({row_reg, col_reg}<18'b001101110010111000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001101110010111000) && ({row_reg, col_reg}<18'b001101110010111110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001101110010111110) && ({row_reg, col_reg}<18'b001101110011000000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001101110011000000) && ({row_reg, col_reg}<18'b001101110011000010)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001101110011000010)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}==18'b001101110011000011)) color_data = 12'b100010111101;
		if(({row_reg, col_reg}==18'b001101110011000100)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==18'b001101110011000101)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b001101110011000110)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}>=18'b001101110011000111) && ({row_reg, col_reg}<18'b001101110011001001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001101110011001001) && ({row_reg, col_reg}<18'b001101110011010010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b001101110011010010) && ({row_reg, col_reg}<18'b001101110011011010)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}>=18'b001101110011011010) && ({row_reg, col_reg}<18'b001101110011011100)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b001101110011011100)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}==18'b001101110011011101)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}>=18'b001101110011011110) && ({row_reg, col_reg}<18'b001101110011100000)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}>=18'b001101110011100000) && ({row_reg, col_reg}<18'b001101110011100100)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b001101110011100100) && ({row_reg, col_reg}<18'b001101111001000110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001101111001000110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001101111001000111) && ({row_reg, col_reg}<18'b001101111001001010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001101111001001010)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001101111001001011)) color_data = 12'b100010111101;
		if(({row_reg, col_reg}==18'b001101111001001100)) color_data = 12'b100110111100;
		if(({row_reg, col_reg}==18'b001101111001001101)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b001101111001001110)) color_data = 12'b101010111011;
		if(({row_reg, col_reg}==18'b001101111001001111)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}==18'b001101111001010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001101111001010001)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}==18'b001101111001010010)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b001101111001010011) && ({row_reg, col_reg}<18'b001101111001101100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001101111001101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001101111001101101) && ({row_reg, col_reg}<18'b001101111010001001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001101111010001001)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b001101111010001010) && ({row_reg, col_reg}<18'b001101111010101110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001101111010101110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b001101111010101111)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001101111010110000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001101111010110001) && ({row_reg, col_reg}<18'b001101111010110011)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b001101111010110011)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==18'b001101111010110100)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b001101111010110101)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b001101111010110110) && ({row_reg, col_reg}<18'b001101111010111000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001101111010111000) && ({row_reg, col_reg}<18'b001101111010111110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001101111010111110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001101111010111111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001101111011000000) && ({row_reg, col_reg}<18'b001101111011000010)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001101111011000010)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}==18'b001101111011000011)) color_data = 12'b100110111101;
		if(({row_reg, col_reg}==18'b001101111011000100)) color_data = 12'b100110111100;
		if(({row_reg, col_reg}>=18'b001101111011000101) && ({row_reg, col_reg}<18'b001101111011000111)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}>=18'b001101111011000111) && ({row_reg, col_reg}<18'b001101111011001101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b001101111011001101) && ({row_reg, col_reg}<18'b001101111011010000)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==18'b001101111011010000)) color_data = 12'b101110011010;
		if(({row_reg, col_reg}>=18'b001101111011010001) && ({row_reg, col_reg}<18'b001101111011010011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001101111011010011) && ({row_reg, col_reg}<18'b001101111011011010)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==18'b001101111011011010)) color_data = 12'b100110011011;
		if(({row_reg, col_reg}==18'b001101111011011011)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b001101111011011100)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}>=18'b001101111011011101) && ({row_reg, col_reg}<18'b001101111011011111)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b001101111011011111)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}>=18'b001101111011100000) && ({row_reg, col_reg}<18'b001101111011100100)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b001101111011100100) && ({row_reg, col_reg}<18'b001110000000110000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001110000000110000)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}>=18'b001110000000110001) && ({row_reg, col_reg}<18'b001110000000110100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001110000000110100) && ({row_reg, col_reg}<18'b001110000000110111)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001110000000110111)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}>=18'b001110000000111000) && ({row_reg, col_reg}<18'b001110000000111010)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b001110000000111010) && ({row_reg, col_reg}<18'b001110000000111110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001110000000111110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001110000000111111)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}>=18'b001110000001000000) && ({row_reg, col_reg}<18'b001110000001000010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001110000001000010) && ({row_reg, col_reg}<18'b001110000001000100)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b001110000001000100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001110000001000101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001110000001000110) && ({row_reg, col_reg}<18'b001110000001001001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001110000001001001)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001110000001001010)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001110000001001011)) color_data = 12'b100110111100;
		if(({row_reg, col_reg}==18'b001110000001001100)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b001110000001001101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001110000001001110)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==18'b001110000001001111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b001110000001010000)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b001110000001010001) && ({row_reg, col_reg}<18'b001110000001101100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001110000001101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001110000001101101) && ({row_reg, col_reg}<18'b001110000010001001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b001110000010001001) && ({row_reg, col_reg}<18'b001110000010101110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001110000010101110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b001110000010101111)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001110000010110000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001110000010110001)) color_data = 12'b101010111010;
		if(({row_reg, col_reg}==18'b001110000010110010)) color_data = 12'b101010111011;
		if(({row_reg, col_reg}==18'b001110000010110011)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b001110000010110100)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b001110000010110101)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b001110000010110110) && ({row_reg, col_reg}<18'b001110000010111000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001110000010111000) && ({row_reg, col_reg}<18'b001110000010111110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001110000010111110) && ({row_reg, col_reg}<18'b001110000011000000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001110000011000000)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}==18'b001110000011000001)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}>=18'b001110000011000010) && ({row_reg, col_reg}<18'b001110000011000100)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==18'b001110000011000100)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b001110000011000101)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}>=18'b001110000011000110) && ({row_reg, col_reg}<18'b001110000011001101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001110000011001101)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}>=18'b001110000011001110) && ({row_reg, col_reg}<18'b001110000011010000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001110000011010000)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b001110000011010001) && ({row_reg, col_reg}<18'b001110000011010111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001110000011010111) && ({row_reg, col_reg}<18'b001110000011011010)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001110000011011010)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001110000011011011)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}>=18'b001110000011011100) && ({row_reg, col_reg}<18'b001110000011011110)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==18'b001110000011011110)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b001110000011011111)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}==18'b001110000011100000)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}>=18'b001110000011100001) && ({row_reg, col_reg}<18'b001110000011100011)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b001110000011100011) && ({row_reg, col_reg}<18'b001110000011100110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001110000011100110) && ({row_reg, col_reg}<18'b001110000011101000)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b001110000011101000) && ({row_reg, col_reg}<18'b001110000011101110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001110000011101110) && ({row_reg, col_reg}<18'b001110000011110000)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b001110000011110000) && ({row_reg, col_reg}<18'b001110001000110100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001110001000110100) && ({row_reg, col_reg}<18'b001110001000111001)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001110001000111001) && ({row_reg, col_reg}<18'b001110001000111100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001110001000111100)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001110001000111101) && ({row_reg, col_reg}<18'b001110001001000010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001110001001000010)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b001110001001000011)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}==18'b001110001001000100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001110001001000101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001110001001000110) && ({row_reg, col_reg}<18'b001110001001001000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001110001001001000) && ({row_reg, col_reg}<18'b001110001001001010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001110001001001010)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001110001001001011)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==18'b001110001001001100)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b001110001001001101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001110001001001110)) color_data = 12'b101010111010;
		if(({row_reg, col_reg}==18'b001110001001001111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b001110001001010000)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b001110001001010001) && ({row_reg, col_reg}<18'b001110001001101100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001110001001101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001110001001101101) && ({row_reg, col_reg}<18'b001110001010001001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001110001010001001)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b001110001010001010) && ({row_reg, col_reg}<18'b001110001010010111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001110001010010111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b001110001010011000) && ({row_reg, col_reg}<18'b001110001010101110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001110001010101110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b001110001010101111)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001110001010110000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001110001010110001)) color_data = 12'b101010111010;
		if(({row_reg, col_reg}==18'b001110001010110010)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b001110001010110011)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b001110001010110100)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b001110001010110101)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b001110001010110110) && ({row_reg, col_reg}<18'b001110001010111000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001110001010111000) && ({row_reg, col_reg}<18'b001110001010111110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001110001010111110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001110001010111111)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b001110001011000000) && ({row_reg, col_reg}<18'b001110001011000010)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b001110001011000010)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==18'b001110001011000011)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b001110001011000100)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b001110001011000101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001110001011000110) && ({row_reg, col_reg}<18'b001110001011001100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001110001011001100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001110001011001101) && ({row_reg, col_reg}<18'b001110001011001111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001110001011001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001110001011010000) && ({row_reg, col_reg}<18'b001110001011010100)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001110001011010100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001110001011010101) && ({row_reg, col_reg}<18'b001110001011011011)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001110001011011011)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}>=18'b001110001011011100) && ({row_reg, col_reg}<18'b001110001011011110)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}==18'b001110001011011110)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==18'b001110001011011111)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}>=18'b001110001011100000) && ({row_reg, col_reg}<18'b001110001011100010)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}>=18'b001110001011100010) && ({row_reg, col_reg}<18'b001110001011100100)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b001110001011100100) && ({row_reg, col_reg}<18'b001110001011100110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001110001011100110) && ({row_reg, col_reg}<18'b001110001011101000)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b001110001011101000) && ({row_reg, col_reg}<18'b001110001011101111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001110001011101111)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b001110001011110000) && ({row_reg, col_reg}<18'b001110010000101110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001110010000101110) && ({row_reg, col_reg}<18'b001110010000110000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001110010000110000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001110010000110001)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001110010000110010) && ({row_reg, col_reg}<18'b001110010000110100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001110010000110100) && ({row_reg, col_reg}<18'b001110010000111011)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001110010000111011)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}==18'b001110010000111100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001110010000111101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001110010000111110) && ({row_reg, col_reg}<18'b001110010001000010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001110010001000010) && ({row_reg, col_reg}<18'b001110010001000100)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b001110010001000100)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}>=18'b001110010001000101) && ({row_reg, col_reg}<18'b001110010001000111)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001110010001000111) && ({row_reg, col_reg}<18'b001110010001001001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001110010001001001)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001110010001001010)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}==18'b001110010001001011)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==18'b001110010001001100)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b001110010001001101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001110010001001110)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==18'b001110010001001111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b001110010001010000)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b001110010001010001) && ({row_reg, col_reg}<18'b001110010001101101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b001110010001101101) && ({row_reg, col_reg}<18'b001110010001101111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b001110010001101111) && ({row_reg, col_reg}<18'b001110010001110001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001110010001110001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001110010001110010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001110010001110011) && ({row_reg, col_reg}<18'b001110010010001001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001110010010001001)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b001110010010001010) && ({row_reg, col_reg}<18'b001110010010101110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001110010010101110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b001110010010101111)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001110010010110000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001110010010110001)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001110010010110010)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b001110010010110011)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b001110010010110100)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b001110010010110101)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001110010010110110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001110010010110111)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}==18'b001110010010111000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001110010010111001) && ({row_reg, col_reg}<18'b001110010010111011)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001110010010111011) && ({row_reg, col_reg}<18'b001110010010111110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001110010010111110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001110010010111111)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b001110010011000000) && ({row_reg, col_reg}<18'b001110010011000010)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b001110010011000010)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==18'b001110010011000011)) color_data = 12'b101010101100;
		if(({row_reg, col_reg}==18'b001110010011000100)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b001110010011000101)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==18'b001110010011000110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001110010011000111)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}>=18'b001110010011001000) && ({row_reg, col_reg}<18'b001110010011001010)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001110010011001010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001110010011001011)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001110010011001100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b001110010011001101) && ({row_reg, col_reg}<18'b001110010011001111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001110010011001111) && ({row_reg, col_reg}<18'b001110010011010001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b001110010011010001)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b001110010011010010) && ({row_reg, col_reg}<18'b001110010011010101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001110010011010101) && ({row_reg, col_reg}<18'b001110010011011001)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001110010011011001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001110010011011010)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001110010011011011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001110010011011100)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==18'b001110010011011101)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}>=18'b001110010011011110) && ({row_reg, col_reg}<18'b001110010011100000)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}>=18'b001110010011100000) && ({row_reg, col_reg}<18'b001110010011100010)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b001110010011100010)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}==18'b001110010011100011)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b001110010011100100) && ({row_reg, col_reg}<18'b001110010011100111)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b001110010011100111) && ({row_reg, col_reg}<18'b001110011000101100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001110011000101100) && ({row_reg, col_reg}<18'b001110011000110010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001110011000110010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001110011000110011) && ({row_reg, col_reg}<18'b001110011000110101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001110011000110101) && ({row_reg, col_reg}<18'b001110011000110111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001110011000110111) && ({row_reg, col_reg}<18'b001110011000111011)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001110011000111011) && ({row_reg, col_reg}<18'b001110011001000010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001110011001000010)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b001110011001000011) && ({row_reg, col_reg}<18'b001110011001001001)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}==18'b001110011001001001)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001110011001001010)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}==18'b001110011001001011)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==18'b001110011001001100)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b001110011001001101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001110011001001110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001110011001001111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001110011001010000)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b001110011001010001) && ({row_reg, col_reg}<18'b001110011001110000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001110011001110000)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==18'b001110011001110001)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001110011001110010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b001110011001110011) && ({row_reg, col_reg}<18'b001110011001110110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b001110011001110110) && ({row_reg, col_reg}<18'b001110011010001000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001110011010001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001110011010001001) && ({row_reg, col_reg}<18'b001110011010101110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001110011010101110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b001110011010101111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001110011010110000) && ({row_reg, col_reg}<18'b001110011010110010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001110011010110010)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b001110011010110011)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b001110011010110100)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}==18'b001110011010110101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001110011010110110) && ({row_reg, col_reg}<18'b001110011010111000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001110011010111000)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b001110011010111001) && ({row_reg, col_reg}<18'b001110011010111110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001110011010111110)) color_data = 12'b011110111110;
		if(({row_reg, col_reg}==18'b001110011010111111)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001110011011000000)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}==18'b001110011011000001)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b001110011011000010)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==18'b001110011011000011)) color_data = 12'b101010111100;
		if(({row_reg, col_reg}==18'b001110011011000100)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b001110011011000101)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==18'b001110011011000110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b001110011011000111) && ({row_reg, col_reg}<18'b001110011011001011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001110011011001011)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==18'b001110011011001100)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b001110011011001101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001110011011001110)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b001110011011001111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001110011011010000)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==18'b001110011011010001)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b001110011011010010) && ({row_reg, col_reg}<18'b001110011011010101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001110011011010101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001110011011010110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001110011011010111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001110011011011000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001110011011011001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001110011011011010) && ({row_reg, col_reg}<18'b001110011011011100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001110011011011100)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==18'b001110011011011101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001110011011011110) && ({row_reg, col_reg}<18'b001110011011100000)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==18'b001110011011100000)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}>=18'b001110011011100001) && ({row_reg, col_reg}<18'b001110011011100011)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}>=18'b001110011011100011) && ({row_reg, col_reg}<18'b001110011011100101)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}>=18'b001110011011100101) && ({row_reg, col_reg}<18'b001110011011100111)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b001110011011100111) && ({row_reg, col_reg}<18'b001110100000101011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001110100000101011) && ({row_reg, col_reg}<18'b001110100000110000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001110100000110000) && ({row_reg, col_reg}<18'b001110100000110010)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}>=18'b001110100000110010) && ({row_reg, col_reg}<18'b001110100000110101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001110100000110101) && ({row_reg, col_reg}<18'b001110100001000010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001110100001000010)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}>=18'b001110100001000011) && ({row_reg, col_reg}<18'b001110100001000101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001110100001000101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001110100001000110) && ({row_reg, col_reg}<18'b001110100001001001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001110100001001001)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001110100001001010)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}==18'b001110100001001011)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==18'b001110100001001100)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b001110100001001101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001110100001001110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001110100001001111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001110100001010000)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b001110100001010001) && ({row_reg, col_reg}<18'b001110100001110001)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001110100001110001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b001110100001110010) && ({row_reg, col_reg}<18'b001110100001110110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b001110100001110110) && ({row_reg, col_reg}<18'b001110100001111011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b001110100001111011) && ({row_reg, col_reg}<18'b001110100001111101)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b001110100001111101) && ({row_reg, col_reg}<18'b001110100010001000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001110100010001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001110100010001001) && ({row_reg, col_reg}<18'b001110100010011011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001110100010011011)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b001110100010011100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001110100010011101) && ({row_reg, col_reg}<18'b001110100010011111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001110100010011111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b001110100010100000) && ({row_reg, col_reg}<18'b001110100010100010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001110100010100010)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b001110100010100011) && ({row_reg, col_reg}<18'b001110100010101011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b001110100010101011) && ({row_reg, col_reg}<18'b001110100010101110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b001110100010101110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b001110100010101111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001110100010110000) && ({row_reg, col_reg}<18'b001110100010110010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001110100010110010)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b001110100010110011)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b001110100010110100)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b001110100010110101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001110100010110110) && ({row_reg, col_reg}<18'b001110100010111001)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b001110100010111001) && ({row_reg, col_reg}<18'b001110100010111110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001110100010111110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001110100010111111)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b001110100011000000) && ({row_reg, col_reg}<18'b001110100011000010)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}==18'b001110100011000010)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}>=18'b001110100011000011) && ({row_reg, col_reg}<18'b001110100011000101)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b001110100011000101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001110100011000110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b001110100011000111) && ({row_reg, col_reg}<18'b001110100011001011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001110100011001011)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b001110100011001100) && ({row_reg, col_reg}<18'b001110100011001110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001110100011001110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001110100011001111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001110100011010000)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==18'b001110100011010001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001110100011010010) && ({row_reg, col_reg}<18'b001110100011010100)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b001110100011010100) && ({row_reg, col_reg}<18'b001110100011010110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001110100011010110)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==18'b001110100011010111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001110100011011000) && ({row_reg, col_reg}<18'b001110100011011010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b001110100011011010) && ({row_reg, col_reg}<18'b001110100011011101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001110100011011101) && ({row_reg, col_reg}<18'b001110100011011111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001110100011011111)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}>=18'b001110100011100000) && ({row_reg, col_reg}<18'b001110100011100011)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b001110100011100011)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b001110100011100100)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}==18'b001110100011100101)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b001110100011100110) && ({row_reg, col_reg}<18'b001110100011101000)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b001110100011101000) && ({row_reg, col_reg}<18'b001110101000101011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001110101000101011) && ({row_reg, col_reg}<18'b001110101000110000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001110101000110000) && ({row_reg, col_reg}<18'b001110101000110010)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}==18'b001110101000110010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001110101000110011) && ({row_reg, col_reg}<18'b001110101000111001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001110101000111001)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b001110101000111010)) color_data = 12'b011110111111;
		if(({row_reg, col_reg}==18'b001110101000111011)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}>=18'b001110101000111100) && ({row_reg, col_reg}<18'b001110101000111110)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b001110101000111110) && ({row_reg, col_reg}<18'b001110101001000000)) color_data = 12'b011110111111;
		if(({row_reg, col_reg}>=18'b001110101001000000) && ({row_reg, col_reg}<18'b001110101001000100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001110101001000100) && ({row_reg, col_reg}<18'b001110101001001001)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==18'b001110101001001001)) color_data = 12'b011110111101;
		if(({row_reg, col_reg}==18'b001110101001001010)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}==18'b001110101001001011)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b001110101001001100)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b001110101001001101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001110101001001110)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==18'b001110101001001111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b001110101001010000)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b001110101001010001) && ({row_reg, col_reg}<18'b001110101001110000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001110101001110000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b001110101001110001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001110101001110010) && ({row_reg, col_reg}<18'b001110101001110110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b001110101001110110) && ({row_reg, col_reg}<18'b001110101010000110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b001110101010000110) && ({row_reg, col_reg}<18'b001110101010001000)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b001110101010001000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001110101010001001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001110101010001010) && ({row_reg, col_reg}<18'b001110101010011011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001110101010011011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b001110101010011100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b001110101010011101) && ({row_reg, col_reg}<18'b001110101010011111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b001110101010011111) && ({row_reg, col_reg}<18'b001110101010101011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b001110101010101011) && ({row_reg, col_reg}<18'b001110101010101110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b001110101010101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001110101010101111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001110101010110000) && ({row_reg, col_reg}<18'b001110101010110010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001110101010110010)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b001110101010110011)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==18'b001110101010110100)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}==18'b001110101010110101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001110101010110110) && ({row_reg, col_reg}<18'b001110101010111000)) color_data = 12'b011010111111;
		if(({row_reg, col_reg}==18'b001110101010111000)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b001110101010111001)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}>=18'b001110101010111010) && ({row_reg, col_reg}<18'b001110101010111110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001110101010111110)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001110101010111111)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}>=18'b001110101011000000) && ({row_reg, col_reg}<18'b001110101011000010)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}==18'b001110101011000010)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}>=18'b001110101011000011) && ({row_reg, col_reg}<18'b001110101011000101)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}>=18'b001110101011000101) && ({row_reg, col_reg}<18'b001110101011000111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b001110101011000111) && ({row_reg, col_reg}<18'b001110101011001001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001110101011001001) && ({row_reg, col_reg}<18'b001110101011001011)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001110101011001011)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}>=18'b001110101011001100) && ({row_reg, col_reg}<18'b001110101011001110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001110101011001110)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b001110101011001111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001110101011010000)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==18'b001110101011010001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001110101011010010) && ({row_reg, col_reg}<18'b001110101011010101)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001110101011010101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001110101011010110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b001110101011010111) && ({row_reg, col_reg}<18'b001110101011011001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001110101011011001)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b001110101011011010) && ({row_reg, col_reg}<18'b001110101011100000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001110101011100000)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==18'b001110101011100001)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}>=18'b001110101011100010) && ({row_reg, col_reg}<18'b001110101011100100)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b001110101011100100)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b001110101011100101)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}==18'b001110101011100110)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001110101011100111)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b001110101011101000) && ({row_reg, col_reg}<18'b001110110000101100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001110110000101100) && ({row_reg, col_reg}<18'b001110110000110000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001110110000110000)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}>=18'b001110110000110001) && ({row_reg, col_reg}<18'b001110110000110101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001110110000110101) && ({row_reg, col_reg}<18'b001110110000111000)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b001110110000111000)) color_data = 12'b010110101110;
		if(({row_reg, col_reg}==18'b001110110000111001)) color_data = 12'b010110101111;
		if(({row_reg, col_reg}>=18'b001110110000111010) && ({row_reg, col_reg}<18'b001110110000111100)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b001110110000111100)) color_data = 12'b011010011111;
		if(({row_reg, col_reg}>=18'b001110110000111101) && ({row_reg, col_reg}<18'b001110110001000000)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b001110110001000000)) color_data = 12'b011010011101;
		if(({row_reg, col_reg}==18'b001110110001000001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001110110001000010)) color_data = 12'b011110111110;
		if(({row_reg, col_reg}==18'b001110110001000011)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}==18'b001110110001000100)) color_data = 12'b010110111100;
		if(({row_reg, col_reg}>=18'b001110110001000101) && ({row_reg, col_reg}<18'b001110110001001001)) color_data = 12'b010110111101;
		if(({row_reg, col_reg}==18'b001110110001001001)) color_data = 12'b011010101100;
		if(({row_reg, col_reg}==18'b001110110001001010)) color_data = 12'b011110101011;
		if(({row_reg, col_reg}==18'b001110110001001011)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b001110110001001100)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b001110110001001101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001110110001001110)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==18'b001110110001001111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b001110110001010000)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b001110110001010001) && ({row_reg, col_reg}<18'b001110110001110000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001110110001110000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b001110110001110001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b001110110001110010) && ({row_reg, col_reg}<18'b001110110001110110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001110110001110110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001110110001110111) && ({row_reg, col_reg}<18'b001110110001111101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b001110110001111101) && ({row_reg, col_reg}<18'b001110110001111111)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b001110110001111111) && ({row_reg, col_reg}<18'b001110110010001000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b001110110010001000) && ({row_reg, col_reg}<18'b001110110010001010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001110110010001010) && ({row_reg, col_reg}<18'b001110110010011100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b001110110010011100) && ({row_reg, col_reg}<18'b001110110010011111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b001110110010011111) && ({row_reg, col_reg}<18'b001110110010100001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001110110010100001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b001110110010100010) && ({row_reg, col_reg}<18'b001110110010101011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b001110110010101011) && ({row_reg, col_reg}<18'b001110110010101110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b001110110010101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001110110010101111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001110110010110000) && ({row_reg, col_reg}<18'b001110110010110010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001110110010110010)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==18'b001110110010110011)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==18'b001110110010110100)) color_data = 12'b011110011100;
		if(({row_reg, col_reg}==18'b001110110010110101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001110110010110110) && ({row_reg, col_reg}<18'b001110110010111000)) color_data = 12'b010110101111;
		if(({row_reg, col_reg}==18'b001110110010111000)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b001110110010111001)) color_data = 12'b011110111111;
		if(({row_reg, col_reg}==18'b001110110010111010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001110110010111011) && ({row_reg, col_reg}<18'b001110110010111101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001110110010111101) && ({row_reg, col_reg}<18'b001110110010111111)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001110110010111111)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}>=18'b001110110011000000) && ({row_reg, col_reg}<18'b001110110011000010)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}>=18'b001110110011000010) && ({row_reg, col_reg}<18'b001110110011000100)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b001110110011000100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001110110011000101) && ({row_reg, col_reg}<18'b001110110011000111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b001110110011000111) && ({row_reg, col_reg}<18'b001110110011001011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001110110011001011)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b001110110011001100)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b001110110011001101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001110110011001110)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b001110110011001111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001110110011010000)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b001110110011010001) && ({row_reg, col_reg}<18'b001110110011010101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b001110110011010101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001110110011010110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b001110110011010111) && ({row_reg, col_reg}<18'b001110110011011001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001110110011011001)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001110110011011010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001110110011011011)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b001110110011011100) && ({row_reg, col_reg}<18'b001110110011100000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001110110011100000) && ({row_reg, col_reg}<18'b001110110011100010)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==18'b001110110011100010)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==18'b001110110011100011)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b001110110011100100)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}==18'b001110110011100101)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b001110110011100110)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}==18'b001110110011100111)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001110110011101000)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b001110110011101001) && ({row_reg, col_reg}<18'b001110111000101110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001110111000101110) && ({row_reg, col_reg}<18'b001110111000110000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001110111000110000) && ({row_reg, col_reg}<18'b001110111000110100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001110111000110100) && ({row_reg, col_reg}<18'b001110111000110111)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b001110111000110111)) color_data = 12'b010110101111;
		if(({row_reg, col_reg}==18'b001110111000111000)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}==18'b001110111000111001)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b001110111000111010)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}>=18'b001110111000111011) && ({row_reg, col_reg}<18'b001110111000111110)) color_data = 12'b010010001110;
		if(({row_reg, col_reg}==18'b001110111000111110)) color_data = 12'b010001111101;
		if(({row_reg, col_reg}==18'b001110111000111111)) color_data = 12'b010001111100;
		if(({row_reg, col_reg}==18'b001110111001000000)) color_data = 12'b010010001011;
		if(({row_reg, col_reg}==18'b001110111001000001)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==18'b001110111001000010)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}>=18'b001110111001000011) && ({row_reg, col_reg}<18'b001110111001001001)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b001110111001001001)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b001110111001001010)) color_data = 12'b101011011110;
		if(({row_reg, col_reg}==18'b001110111001001011)) color_data = 12'b100110111011;
		if(({row_reg, col_reg}>=18'b001110111001001100) && ({row_reg, col_reg}<18'b001110111001001110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001110111001001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==18'b001110111001001111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b001110111001010000)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b001110111001010001) && ({row_reg, col_reg}<18'b001110111001101011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001110111001101011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b001110111001101100) && ({row_reg, col_reg}<18'b001110111001101110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001110111001101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001110111001101111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001110111001110000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001110111001110001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b001110111001110010) && ({row_reg, col_reg}<18'b001110111001110101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001110111001110101) && ({row_reg, col_reg}<18'b001110111001111000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001110111001111000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001110111001111001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001110111001111010) && ({row_reg, col_reg}<18'b001110111001111110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001110111001111110)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==18'b001110111001111111)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b001110111010000000) && ({row_reg, col_reg}<18'b001110111010000100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001110111010000100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b001110111010000101) && ({row_reg, col_reg}<18'b001110111010010010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001110111010010010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001110111010010011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b001110111010010100) && ({row_reg, col_reg}<18'b001110111010010110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001110111010010110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b001110111010010111) && ({row_reg, col_reg}<18'b001110111010011010)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001110111010011010) && ({row_reg, col_reg}<18'b001110111010011101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b001110111010011101) && ({row_reg, col_reg}<18'b001110111010011111)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==18'b001110111010011111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b001110111010100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b001110111010100001) && ({row_reg, col_reg}<18'b001110111010101101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001110111010101101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b001110111010101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001110111010101111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001110111010110000) && ({row_reg, col_reg}<18'b001110111010110010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001110111010110010)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b001110111010110011)) color_data = 12'b100010011011;
		if(({row_reg, col_reg}==18'b001110111010110100)) color_data = 12'b010110001011;
		if(({row_reg, col_reg}==18'b001110111010110101)) color_data = 12'b010010001100;
		if(({row_reg, col_reg}>=18'b001110111010110110) && ({row_reg, col_reg}<18'b001110111010111000)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b001110111010111000)) color_data = 12'b010010011110;
		if(({row_reg, col_reg}==18'b001110111010111001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001110111010111010) && ({row_reg, col_reg}<18'b001110111010111100)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}==18'b001110111010111100)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b001110111010111101) && ({row_reg, col_reg}<18'b001110111010111111)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}==18'b001110111010111111)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}>=18'b001110111011000000) && ({row_reg, col_reg}<18'b001110111011000011)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}>=18'b001110111011000011) && ({row_reg, col_reg}<18'b001110111011000110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001110111011000110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001110111011000111)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b001110111011001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b001110111011001001)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b001110111011001010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b001110111011001011)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b001110111011001100) && ({row_reg, col_reg}<18'b001110111011001110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001110111011001110) && ({row_reg, col_reg}<18'b001110111011010001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b001110111011010001) && ({row_reg, col_reg}<18'b001110111011010100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b001110111011010100)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b001110111011010101)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b001110111011010110) && ({row_reg, col_reg}<18'b001110111011011010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b001110111011011010) && ({row_reg, col_reg}<18'b001110111011011100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001110111011011100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b001110111011011101) && ({row_reg, col_reg}<18'b001110111011011111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001110111011011111) && ({row_reg, col_reg}<18'b001110111011100010)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001110111011100010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001110111011100011) && ({row_reg, col_reg}<18'b001110111011100101)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==18'b001110111011100101)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}>=18'b001110111011100110) && ({row_reg, col_reg}<18'b001110111011101000)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b001110111011101000)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b001110111011101001) && ({row_reg, col_reg}<18'b001110111011101011)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b001110111011101011) && ({row_reg, col_reg}<18'b001111000000110101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001111000000110101)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b001111000000110110)) color_data = 12'b011010111111;
		if(({row_reg, col_reg}==18'b001111000000110111)) color_data = 12'b010110101111;
		if(({row_reg, col_reg}==18'b001111000000111000)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b001111000000111001)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b001111000000111010) && ({row_reg, col_reg}<18'b001111000000111111)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b001111000000111111)) color_data = 12'b001001101011;
		if(({row_reg, col_reg}==18'b001111000001000000)) color_data = 12'b001001111010;
		if(({row_reg, col_reg}==18'b001111000001000001)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==18'b001111000001000010)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b001111000001000011) && ({row_reg, col_reg}<18'b001111000001001001)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b001111000001001001)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b001111000001001010)) color_data = 12'b101011101110;
		if(({row_reg, col_reg}==18'b001111000001001011)) color_data = 12'b100110111011;
		if(({row_reg, col_reg}==18'b001111000001001100)) color_data = 12'b101010111010;
		if(({row_reg, col_reg}==18'b001111000001001101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001111000001001110)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==18'b001111000001001111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b001111000001010000)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b001111000001010001) && ({row_reg, col_reg}<18'b001111000001101110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001111000001101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001111000001101111) && ({row_reg, col_reg}<18'b001111000001110001)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001111000001110001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001111000001110010) && ({row_reg, col_reg}<18'b001111000001110111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001111000001110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001111000001111000) && ({row_reg, col_reg}<18'b001111000001111010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b001111000001111010) && ({row_reg, col_reg}<18'b001111000001111100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001111000001111100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001111000001111101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001111000001111110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001111000001111111)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b001111000010000000) && ({row_reg, col_reg}<18'b001111000010000100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b001111000010000100) && ({row_reg, col_reg}<18'b001111000010001111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001111000010001111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b001111000010010000) && ({row_reg, col_reg}<18'b001111000010010010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001111000010010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b001111000010010011) && ({row_reg, col_reg}<18'b001111000010011011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001111000010011011)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001111000010011100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001111000010011101)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b001111000010011110) && ({row_reg, col_reg}<18'b001111000010100000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001111000010100000)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b001111000010100001)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b001111000010100010) && ({row_reg, col_reg}<18'b001111000010101101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001111000010101101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b001111000010101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001111000010101111) && ({row_reg, col_reg}<18'b001111000010110001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001111000010110001)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==18'b001111000010110010)) color_data = 12'b101010101100;
		if(({row_reg, col_reg}==18'b001111000010110011)) color_data = 12'b100110011100;
		if(({row_reg, col_reg}==18'b001111000010110100)) color_data = 12'b010101111010;
		if(({row_reg, col_reg}>=18'b001111000010110101) && ({row_reg, col_reg}<18'b001111000010110111)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b001111000010110111)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b001111000010111000)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b001111000010111001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001111000010111010) && ({row_reg, col_reg}<18'b001111000010111101)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001111000010111101)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}>=18'b001111000010111110) && ({row_reg, col_reg}<18'b001111000011000000)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}>=18'b001111000011000000) && ({row_reg, col_reg}<18'b001111000011000010)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b001111000011000010)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==18'b001111000011000011)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}>=18'b001111000011000100) && ({row_reg, col_reg}<18'b001111000011000110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001111000011000110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b001111000011000111) && ({row_reg, col_reg}<18'b001111000011001010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b001111000011001010) && ({row_reg, col_reg}<18'b001111000011001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001111000011001100) && ({row_reg, col_reg}<18'b001111000011001110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001111000011001110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001111000011001111) && ({row_reg, col_reg}<18'b001111000011010001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001111000011010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001111000011010010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001111000011010011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001111000011010100)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b001111000011010101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001111000011010110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==18'b001111000011010111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001111000011011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001111000011011001) && ({row_reg, col_reg}<18'b001111000011011110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001111000011011110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001111000011011111) && ({row_reg, col_reg}<18'b001111000011100011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001111000011100011)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==18'b001111000011100100)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==18'b001111000011100101)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b001111000011100110)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}==18'b001111000011100111)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b001111000011101000)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}==18'b001111000011101001)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b001111000011101010) && ({row_reg, col_reg}<18'b001111000011101101)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b001111000011101101) && ({row_reg, col_reg}<18'b001111001000110110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001111001000110110)) color_data = 12'b011110111111;
		if(({row_reg, col_reg}==18'b001111001000110111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001111001000111000)) color_data = 12'b010010001100;
		if(({row_reg, col_reg}==18'b001111001000111001)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}>=18'b001111001000111010) && ({row_reg, col_reg}<18'b001111001000111101)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b001111001000111101) && ({row_reg, col_reg}<18'b001111001000111111)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b001111001000111111)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b001111001001000000)) color_data = 12'b001010001010;
		if(({row_reg, col_reg}==18'b001111001001000001)) color_data = 12'b010110111101;
		if(({row_reg, col_reg}==18'b001111001001000010)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b001111001001000011) && ({row_reg, col_reg}<18'b001111001001001000)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b001111001001001000) && ({row_reg, col_reg}<18'b001111001001001010)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b001111001001001010)) color_data = 12'b101011101111;
		if(({row_reg, col_reg}==18'b001111001001001011)) color_data = 12'b100110111011;
		if(({row_reg, col_reg}>=18'b001111001001001100) && ({row_reg, col_reg}<18'b001111001001001110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001111001001001110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001111001001001111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b001111001001010000) && ({row_reg, col_reg}<18'b001111001001101100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001111001001101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001111001001101101) && ({row_reg, col_reg}<18'b001111001001101111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001111001001101111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b001111001001110000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001111001001110001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001111001001110010) && ({row_reg, col_reg}<18'b001111001001111011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b001111001001111011) && ({row_reg, col_reg}<18'b001111001001111111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001111001001111111)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b001111001010000000) && ({row_reg, col_reg}<18'b001111001010000100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001111001010000100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b001111001010000101) && ({row_reg, col_reg}<18'b001111001010010010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001111001010010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b001111001010010011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001111001010010100)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b001111001010010101) && ({row_reg, col_reg}<18'b001111001010011000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001111001010011000)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b001111001010011001) && ({row_reg, col_reg}<18'b001111001010011110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001111001010011110)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001111001010011111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001111001010100000)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b001111001010100001)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001111001010100010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b001111001010100011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001111001010100100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b001111001010100101) && ({row_reg, col_reg}<18'b001111001010101110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001111001010101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001111001010101111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001111001010110000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001111001010110001)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==18'b001111001010110010)) color_data = 12'b101010101100;
		if(({row_reg, col_reg}==18'b001111001010110011)) color_data = 12'b100110011100;
		if(({row_reg, col_reg}==18'b001111001010110100)) color_data = 12'b010101111011;
		if(({row_reg, col_reg}==18'b001111001010110101)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b001111001010110110)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b001111001010110111)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b001111001010111000)) color_data = 12'b010010011101;
		if(({row_reg, col_reg}==18'b001111001010111001)) color_data = 12'b011110111110;
		if(({row_reg, col_reg}==18'b001111001010111010)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001111001010111011)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}==18'b001111001010111100)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}>=18'b001111001010111101) && ({row_reg, col_reg}<18'b001111001010111111)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}>=18'b001111001010111111) && ({row_reg, col_reg}<18'b001111001011000010)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}>=18'b001111001011000010) && ({row_reg, col_reg}<18'b001111001011000100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001111001011000100) && ({row_reg, col_reg}<18'b001111001011000111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001111001011000111) && ({row_reg, col_reg}<18'b001111001011001100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001111001011001100)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b001111001011001101) && ({row_reg, col_reg}<18'b001111001011010011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001111001011010011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001111001011010100)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b001111001011010101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001111001011010110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==18'b001111001011010111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001111001011011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001111001011011001) && ({row_reg, col_reg}<18'b001111001011011110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001111001011011110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001111001011011111) && ({row_reg, col_reg}<18'b001111001011100001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001111001011100001)) color_data = 12'b101110011001;
		if(({row_reg, col_reg}>=18'b001111001011100010) && ({row_reg, col_reg}<18'b001111001011100100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001111001011100100)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}>=18'b001111001011100101) && ({row_reg, col_reg}<18'b001111001011100111)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==18'b001111001011100111)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}==18'b001111001011101000)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b001111001011101001)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}>=18'b001111001011101010) && ({row_reg, col_reg}<18'b001111001011101100)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001111001011101100)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b001111001011101101) && ({row_reg, col_reg}<18'b001111010000110000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001111010000110000) && ({row_reg, col_reg}<18'b001111010000110100)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001111010000110100)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}==18'b001111010000110101)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001111010000110110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001111010000110111)) color_data = 12'b011010011101;
		if(({row_reg, col_reg}==18'b001111010000111000)) color_data = 12'b010001111011;
		if(({row_reg, col_reg}==18'b001111010000111001)) color_data = 12'b001101101010;
		if(({row_reg, col_reg}>=18'b001111010000111010) && ({row_reg, col_reg}<18'b001111010000111100)) color_data = 12'b001101111011;
		if(({row_reg, col_reg}>=18'b001111010000111100) && ({row_reg, col_reg}<18'b001111010000111111)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b001111010000111111)) color_data = 12'b000101111010;
		if(({row_reg, col_reg}==18'b001111010001000000)) color_data = 12'b000110001010;
		if(({row_reg, col_reg}==18'b001111010001000001)) color_data = 12'b010110111110;
		if(({row_reg, col_reg}==18'b001111010001000010)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b001111010001000011) && ({row_reg, col_reg}<18'b001111010001000101)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b001111010001000101) && ({row_reg, col_reg}<18'b001111010001000111)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b001111010001000111)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b001111010001001000) && ({row_reg, col_reg}<18'b001111010001001010)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b001111010001001010)) color_data = 12'b101011101111;
		if(({row_reg, col_reg}==18'b001111010001001011)) color_data = 12'b100110111100;
		if(({row_reg, col_reg}==18'b001111010001001100)) color_data = 12'b101010111011;
		if(({row_reg, col_reg}==18'b001111010001001101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001111010001001110)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==18'b001111010001001111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b001111010001010000) && ({row_reg, col_reg}<18'b001111010001101011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001111010001101011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b001111010001101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001111010001101101) && ({row_reg, col_reg}<18'b001111010001110000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001111010001110000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001111010001110001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001111010001110010) && ({row_reg, col_reg}<18'b001111010001110110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001111010001110110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001111010001110111) && ({row_reg, col_reg}<18'b001111010001111011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b001111010001111011) && ({row_reg, col_reg}<18'b001111010001111111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001111010001111111)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b001111010010000000) && ({row_reg, col_reg}<18'b001111010010000010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001111010010000010) && ({row_reg, col_reg}<18'b001111010010000100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b001111010010000100) && ({row_reg, col_reg}<18'b001111010010010000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001111010010010000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b001111010010010001)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001111010010010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b001111010010010011) && ({row_reg, col_reg}<18'b001111010010011011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001111010010011011)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b001111010010011100) && ({row_reg, col_reg}<18'b001111010010011110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001111010010011110) && ({row_reg, col_reg}<18'b001111010010100000)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001111010010100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b001111010010100001)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001111010010100010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b001111010010100011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001111010010100100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b001111010010100101) && ({row_reg, col_reg}<18'b001111010010101110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001111010010101110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b001111010010101111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001111010010110000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001111010010110001)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==18'b001111010010110010)) color_data = 12'b101010101100;
		if(({row_reg, col_reg}==18'b001111010010110011)) color_data = 12'b100110011100;
		if(({row_reg, col_reg}==18'b001111010010110100)) color_data = 12'b010101101011;
		if(({row_reg, col_reg}==18'b001111010010110101)) color_data = 12'b010001111100;
		if(({row_reg, col_reg}==18'b001111010010110110)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b001111010010110111)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b001111010010111000)) color_data = 12'b010010001100;
		if(({row_reg, col_reg}==18'b001111010010111001)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001111010010111010)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}>=18'b001111010010111011) && ({row_reg, col_reg}<18'b001111010010111101)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}==18'b001111010010111101)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}>=18'b001111010010111110) && ({row_reg, col_reg}<18'b001111010011000010)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b001111010011000010)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==18'b001111010011000011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001111010011000100) && ({row_reg, col_reg}<18'b001111010011000111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001111010011000111) && ({row_reg, col_reg}<18'b001111010011010100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001111010011010100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b001111010011010101)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b001111010011010110) && ({row_reg, col_reg}<18'b001111010011011000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b001111010011011000) && ({row_reg, col_reg}<18'b001111010011011111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001111010011011111)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b001111010011100000) && ({row_reg, col_reg}<18'b001111010011100010)) color_data = 12'b101110011001;
		if(({row_reg, col_reg}>=18'b001111010011100010) && ({row_reg, col_reg}<18'b001111010011100101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001111010011100101)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==18'b001111010011100110)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}==18'b001111010011100111)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b001111010011101000)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}==18'b001111010011101001)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b001111010011101010)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}>=18'b001111010011101011) && ({row_reg, col_reg}<18'b001111010011101101)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001111010011101101)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b001111010011101110) && ({row_reg, col_reg}<18'b001111011000110000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001111011000110000) && ({row_reg, col_reg}<18'b001111011000110110)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001111011000110110)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}==18'b001111011000110111)) color_data = 12'b011110011100;
		if(({row_reg, col_reg}==18'b001111011000111000)) color_data = 12'b011110011011;
		if(({row_reg, col_reg}>=18'b001111011000111001) && ({row_reg, col_reg}<18'b001111011000111011)) color_data = 12'b011010001011;
		if(({row_reg, col_reg}==18'b001111011000111011)) color_data = 12'b011010011100;
		if(({row_reg, col_reg}==18'b001111011000111100)) color_data = 12'b010010001011;
		if(({row_reg, col_reg}==18'b001111011000111101)) color_data = 12'b010110101101;
		if(({row_reg, col_reg}==18'b001111011000111110)) color_data = 12'b010010101100;
		if(({row_reg, col_reg}==18'b001111011000111111)) color_data = 12'b001110101100;
		if(({row_reg, col_reg}==18'b001111011001000000)) color_data = 12'b010010111110;
		if(({row_reg, col_reg}==18'b001111011001000001)) color_data = 12'b010110111110;
		if(({row_reg, col_reg}>=18'b001111011001000010) && ({row_reg, col_reg}<18'b001111011001000100)) color_data = 12'b011011011111;
		if(({row_reg, col_reg}>=18'b001111011001000100) && ({row_reg, col_reg}<18'b001111011001000110)) color_data = 12'b011011001111;
		if(({row_reg, col_reg}>=18'b001111011001000110) && ({row_reg, col_reg}<18'b001111011001001010)) color_data = 12'b011111001111;
		if(({row_reg, col_reg}==18'b001111011001001010)) color_data = 12'b100011001110;
		if(({row_reg, col_reg}==18'b001111011001001011)) color_data = 12'b100110111100;
		if(({row_reg, col_reg}==18'b001111011001001100)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b001111011001001101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001111011001001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==18'b001111011001001111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b001111011001010000) && ({row_reg, col_reg}<18'b001111011001101000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001111011001101000)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b001111011001101001) && ({row_reg, col_reg}<18'b001111011001101100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001111011001101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b001111011001101101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001111011001101110)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b001111011001101111) && ({row_reg, col_reg}<18'b001111011001110001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b001111011001110001)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b001111011001110010) && ({row_reg, col_reg}<18'b001111011001110101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001111011001110101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001111011001110110) && ({row_reg, col_reg}<18'b001111011001111000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b001111011001111000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001111011001111001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b001111011001111010) && ({row_reg, col_reg}<18'b001111011001111111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001111011001111111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b001111011010000000) && ({row_reg, col_reg}<18'b001111011010000100)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b001111011010000100) && ({row_reg, col_reg}<18'b001111011010001101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001111011010001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001111011010001110) && ({row_reg, col_reg}<18'b001111011010010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b001111011010010000) && ({row_reg, col_reg}<18'b001111011010010010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001111011010010010)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b001111011010010011) && ({row_reg, col_reg}<18'b001111011010010110)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b001111011010010110) && ({row_reg, col_reg}<18'b001111011010011001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001111011010011001) && ({row_reg, col_reg}<18'b001111011010011100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001111011010011100) && ({row_reg, col_reg}<18'b001111011010011111)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001111011010011111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001111011010100000)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==18'b001111011010100001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b001111011010100010) && ({row_reg, col_reg}<18'b001111011010100100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001111011010100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b001111011010100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001111011010100110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b001111011010100111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b001111011010101000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001111011010101001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b001111011010101010) && ({row_reg, col_reg}<18'b001111011010101110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001111011010101110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b001111011010101111)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b001111011010110000) && ({row_reg, col_reg}<18'b001111011010110010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001111011010110010)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b001111011010110011)) color_data = 12'b100110011100;
		if(({row_reg, col_reg}==18'b001111011010110100)) color_data = 12'b010101101011;
		if(({row_reg, col_reg}==18'b001111011010110101)) color_data = 12'b010001111100;
		if(({row_reg, col_reg}==18'b001111011010110110)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b001111011010110111)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b001111011010111000)) color_data = 12'b010110011100;
		if(({row_reg, col_reg}==18'b001111011010111001)) color_data = 12'b100010111101;
		if(({row_reg, col_reg}==18'b001111011010111010)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}>=18'b001111011010111011) && ({row_reg, col_reg}<18'b001111011010111101)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}>=18'b001111011010111101) && ({row_reg, col_reg}<18'b001111011011000000)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b001111011011000000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001111011011000001)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}>=18'b001111011011000010) && ({row_reg, col_reg}<18'b001111011011000100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b001111011011000100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001111011011000101)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==18'b001111011011000110)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b001111011011000111) && ({row_reg, col_reg}<18'b001111011011001011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b001111011011001011) && ({row_reg, col_reg}<18'b001111011011001111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001111011011001111) && ({row_reg, col_reg}<18'b001111011011010010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b001111011011010010) && ({row_reg, col_reg}<18'b001111011011010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001111011011010100)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b001111011011010101)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001111011011010110)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==18'b001111011011010111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b001111011011011000) && ({row_reg, col_reg}<18'b001111011011100000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001111011011100000)) color_data = 12'b101110011001;
		if(({row_reg, col_reg}==18'b001111011011100001)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}>=18'b001111011011100010) && ({row_reg, col_reg}<18'b001111011011100100)) color_data = 12'b101110011001;
		if(({row_reg, col_reg}==18'b001111011011100100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001111011011100101) && ({row_reg, col_reg}<18'b001111011011100111)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==18'b001111011011100111)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}>=18'b001111011011101000) && ({row_reg, col_reg}<18'b001111011011101010)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}>=18'b001111011011101010) && ({row_reg, col_reg}<18'b001111011011101100)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}>=18'b001111011011101100) && ({row_reg, col_reg}<18'b001111011011101110)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001111011011101110)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b001111011011101111) && ({row_reg, col_reg}<18'b001111100000110000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001111100000110000) && ({row_reg, col_reg}<18'b001111100000110011)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b001111100000110011) && ({row_reg, col_reg}<18'b001111100000110110)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}>=18'b001111100000110110) && ({row_reg, col_reg}<18'b001111100000111001)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b001111100000111001)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==18'b001111100000111010)) color_data = 12'b100110111100;
		if(({row_reg, col_reg}==18'b001111100000111011)) color_data = 12'b100110111101;
		if(({row_reg, col_reg}==18'b001111100000111100)) color_data = 12'b100011001101;
		if(({row_reg, col_reg}==18'b001111100000111101)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}>=18'b001111100000111110) && ({row_reg, col_reg}<18'b001111100001000000)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b001111100001000000)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b001111100001000001)) color_data = 12'b010010101101;
		if(({row_reg, col_reg}==18'b001111100001000010)) color_data = 12'b000101111011;
		if(({row_reg, col_reg}>=18'b001111100001000011) && ({row_reg, col_reg}<18'b001111100001000110)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}>=18'b001111100001000110) && ({row_reg, col_reg}<18'b001111100001001001)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b001111100001001001)) color_data = 12'b001110001011;
		if(({row_reg, col_reg}==18'b001111100001001010)) color_data = 12'b010010001010;
		if(({row_reg, col_reg}==18'b001111100001001011)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}==18'b001111100001001100)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b001111100001001101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001111100001001110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==18'b001111100001001111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001111100001010000) && ({row_reg, col_reg}<18'b001111100001101100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001111100001101100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001111100001101101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001111100001101110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001111100001101111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=18'b001111100001110000) && ({row_reg, col_reg}<18'b001111100001110101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001111100001110101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001111100001110110) && ({row_reg, col_reg}<18'b001111100001111000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001111100001111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001111100001111001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b001111100001111010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b001111100001111011) && ({row_reg, col_reg}<18'b001111100010000100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001111100010000100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001111100010000101) && ({row_reg, col_reg}<18'b001111100010001101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001111100010001101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b001111100010001110) && ({row_reg, col_reg}<18'b001111100010010010)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001111100010010010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001111100010010011) && ({row_reg, col_reg}<18'b001111100010011010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b001111100010011010) && ({row_reg, col_reg}<18'b001111100010011100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001111100010011100)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001111100010011101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001111100010011110) && ({row_reg, col_reg}<18'b001111100010100000)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b001111100010100000) && ({row_reg, col_reg}<18'b001111100010100010)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001111100010100010) && ({row_reg, col_reg}<18'b001111100010100100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b001111100010100100)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001111100010100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b001111100010100110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b001111100010100111) && ({row_reg, col_reg}<18'b001111100010101001)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b001111100010101001) && ({row_reg, col_reg}<18'b001111100010101101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b001111100010101101) && ({row_reg, col_reg}<18'b001111100010101111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b001111100010101111) && ({row_reg, col_reg}<18'b001111100010110001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001111100010110001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==18'b001111100010110010)) color_data = 12'b101010101100;
		if(({row_reg, col_reg}==18'b001111100010110011)) color_data = 12'b100110011100;
		if(({row_reg, col_reg}==18'b001111100010110100)) color_data = 12'b010101111011;
		if(({row_reg, col_reg}==18'b001111100010110101)) color_data = 12'b010001111100;
		if(({row_reg, col_reg}==18'b001111100010110110)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b001111100010110111)) color_data = 12'b001101111011;
		if(({row_reg, col_reg}==18'b001111100010111000)) color_data = 12'b011010011100;
		if(({row_reg, col_reg}==18'b001111100010111001)) color_data = 12'b100010111101;
		if(({row_reg, col_reg}==18'b001111100010111010)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==18'b001111100010111011)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b001111100010111100)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b001111100010111101)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}>=18'b001111100010111110) && ({row_reg, col_reg}<18'b001111100011000000)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==18'b001111100011000000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001111100011000001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001111100011000010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b001111100011000011) && ({row_reg, col_reg}<18'b001111100011001011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001111100011001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001111100011001100) && ({row_reg, col_reg}<18'b001111100011010001)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001111100011010001)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b001111100011010010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001111100011010011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b001111100011010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001111100011010101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001111100011010110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001111100011010111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001111100011011000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b001111100011011001) && ({row_reg, col_reg}<18'b001111100011011111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001111100011011111) && ({row_reg, col_reg}<18'b001111100011100010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001111100011100010)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==18'b001111100011100011)) color_data = 12'b101110011001;
		if(({row_reg, col_reg}>=18'b001111100011100100) && ({row_reg, col_reg}<18'b001111100011100111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001111100011100111)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}==18'b001111100011101000)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==18'b001111100011101001)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}>=18'b001111100011101010) && ({row_reg, col_reg}<18'b001111100011101100)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}==18'b001111100011101100)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}>=18'b001111100011101101) && ({row_reg, col_reg}<18'b001111100011110000)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b001111100011110000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001111100011110001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001111100011110010)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b001111100011110011) && ({row_reg, col_reg}<18'b001111101000101111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b001111101000101111)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001111101000110000) && ({row_reg, col_reg}<18'b001111101000110100)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b001111101000110100)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b001111101000110101)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}>=18'b001111101000110110) && ({row_reg, col_reg}<18'b001111101000111001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001111101000111001) && ({row_reg, col_reg}<18'b001111101000111011)) color_data = 12'b101010111011;
		if(({row_reg, col_reg}==18'b001111101000111011)) color_data = 12'b100010111011;
		if(({row_reg, col_reg}==18'b001111101000111100)) color_data = 12'b100111001100;
		if(({row_reg, col_reg}==18'b001111101000111101)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}==18'b001111101000111110)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b001111101000111111)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b001111101001000000)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b001111101001000001)) color_data = 12'b010110111110;
		if(({row_reg, col_reg}==18'b001111101001000010)) color_data = 12'b000110001011;
		if(({row_reg, col_reg}>=18'b001111101001000011) && ({row_reg, col_reg}<18'b001111101001000101)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b001111101001000101)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b001111101001000110)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b001111101001000111) && ({row_reg, col_reg}<18'b001111101001001001)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b001111101001001001)) color_data = 12'b001110001011;
		if(({row_reg, col_reg}==18'b001111101001001010)) color_data = 12'b010001111010;
		if(({row_reg, col_reg}==18'b001111101001001011)) color_data = 12'b100110111100;
		if(({row_reg, col_reg}==18'b001111101001001100)) color_data = 12'b101010111011;
		if(({row_reg, col_reg}==18'b001111101001001101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001111101001001110)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==18'b001111101001001111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b001111101001010000) && ({row_reg, col_reg}<18'b001111101001101100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001111101001101100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001111101001101101) && ({row_reg, col_reg}<18'b001111101001110000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001111101001110000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001111101001110001)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b001111101001110010) && ({row_reg, col_reg}<18'b001111101001110100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001111101001110100)) color_data = 12'b110010111011;
		if(({row_reg, col_reg}==18'b001111101001110101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001111101001110110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001111101001110111) && ({row_reg, col_reg}<18'b001111101001111001)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001111101001111001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b001111101001111010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b001111101001111011) && ({row_reg, col_reg}<18'b001111101001111110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001111101001111110)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001111101001111111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001111101010000000) && ({row_reg, col_reg}<18'b001111101010000010)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001111101010000010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001111101010000011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001111101010000100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b001111101010000101) && ({row_reg, col_reg}<18'b001111101010001101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001111101010001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b001111101010001110) && ({row_reg, col_reg}<18'b001111101010010000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001111101010010000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001111101010010001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001111101010010010) && ({row_reg, col_reg}<18'b001111101010011100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001111101010011100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001111101010011101) && ({row_reg, col_reg}<18'b001111101010011111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001111101010011111)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b001111101010100000) && ({row_reg, col_reg}<18'b001111101010100010)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001111101010100010)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b001111101010100011) && ({row_reg, col_reg}<18'b001111101010100101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001111101010100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b001111101010100110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b001111101010100111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001111101010101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001111101010101001) && ({row_reg, col_reg}<18'b001111101010101101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b001111101010101101) && ({row_reg, col_reg}<18'b001111101010101111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b001111101010101111)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001111101010110000)) color_data = 12'b100110101001;
		if(({row_reg, col_reg}==18'b001111101010110001)) color_data = 12'b101010111010;
		if(({row_reg, col_reg}==18'b001111101010110010)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b001111101010110011)) color_data = 12'b100010011100;
		if(({row_reg, col_reg}==18'b001111101010110100)) color_data = 12'b010001101011;
		if(({row_reg, col_reg}==18'b001111101010110101)) color_data = 12'b010001111100;
		if(({row_reg, col_reg}==18'b001111101010110110)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b001111101010110111)) color_data = 12'b001101111011;
		if(({row_reg, col_reg}==18'b001111101010111000)) color_data = 12'b011010011100;
		if(({row_reg, col_reg}==18'b001111101010111001)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}>=18'b001111101010111010) && ({row_reg, col_reg}<18'b001111101010111101)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}>=18'b001111101010111101) && ({row_reg, col_reg}<18'b001111101010111111)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==18'b001111101010111111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b001111101011000000) && ({row_reg, col_reg}<18'b001111101011000010)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001111101011000010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001111101011000011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001111101011000100) && ({row_reg, col_reg}<18'b001111101011001010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001111101011001010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b001111101011001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001111101011001100) && ({row_reg, col_reg}<18'b001111101011010011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001111101011010011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b001111101011010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001111101011010101)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b001111101011010110) && ({row_reg, col_reg}<18'b001111101011011001)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b001111101011011001) && ({row_reg, col_reg}<18'b001111101011011101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001111101011011101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001111101011011110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001111101011011111) && ({row_reg, col_reg}<18'b001111101011100011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001111101011100011)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b001111101011100100) && ({row_reg, col_reg}<18'b001111101011100111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001111101011100111) && ({row_reg, col_reg}<18'b001111101011101001)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==18'b001111101011101001)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}==18'b001111101011101010)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b001111101011101011)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}>=18'b001111101011101100) && ({row_reg, col_reg}<18'b001111101011101111)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b001111101011101111)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b001111101011110000) && ({row_reg, col_reg}<18'b001111101011110100)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b001111101011110100) && ({row_reg, col_reg}<18'b001111110000101101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001111110000101101) && ({row_reg, col_reg}<18'b001111110000110000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b001111110000110000)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}>=18'b001111110000110001) && ({row_reg, col_reg}<18'b001111110000110011)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}==18'b001111110000110011)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}>=18'b001111110000110100) && ({row_reg, col_reg}<18'b001111110000110110)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}>=18'b001111110000110110) && ({row_reg, col_reg}<18'b001111110000111000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001111110000111000) && ({row_reg, col_reg}<18'b001111110000111011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001111110000111011)) color_data = 12'b100010101001;
		if(({row_reg, col_reg}==18'b001111110000111100)) color_data = 12'b100111001011;
		if(({row_reg, col_reg}==18'b001111110000111101)) color_data = 12'b101111101110;
		if(({row_reg, col_reg}==18'b001111110000111110)) color_data = 12'b101011101110;
		if(({row_reg, col_reg}==18'b001111110000111111)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b001111110001000000)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b001111110001000001)) color_data = 12'b010110111110;
		if(({row_reg, col_reg}==18'b001111110001000010)) color_data = 12'b000101111011;
		if(({row_reg, col_reg}>=18'b001111110001000011) && ({row_reg, col_reg}<18'b001111110001000101)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}>=18'b001111110001000101) && ({row_reg, col_reg}<18'b001111110001001001)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b001111110001001001)) color_data = 12'b001110001011;
		if(({row_reg, col_reg}==18'b001111110001001010)) color_data = 12'b010001111010;
		if(({row_reg, col_reg}==18'b001111110001001011)) color_data = 12'b100110111100;
		if(({row_reg, col_reg}>=18'b001111110001001100) && ({row_reg, col_reg}<18'b001111110001001110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001111110001001110)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==18'b001111110001001111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b001111110001010000) && ({row_reg, col_reg}<18'b001111110001101100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001111110001101100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001111110001101101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b001111110001101110) && ({row_reg, col_reg}<18'b001111110001110000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001111110001110000) && ({row_reg, col_reg}<18'b001111110001110011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001111110001110011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001111110001110100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==18'b001111110001110101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001111110001110110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b001111110001110111) && ({row_reg, col_reg}<18'b001111110001111010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001111110001111010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001111110001111011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001111110001111100) && ({row_reg, col_reg}<18'b001111110010000100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001111110010000100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001111110010000101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001111110010000110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b001111110010000111) && ({row_reg, col_reg}<18'b001111110010001010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001111110010001010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b001111110010001011) && ({row_reg, col_reg}<18'b001111110010001101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001111110010001101)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b001111110010001110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001111110010001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001111110010010000) && ({row_reg, col_reg}<18'b001111110010010011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001111110010010011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001111110010010100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001111110010010101) && ({row_reg, col_reg}<18'b001111110010011100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001111110010011100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001111110010011101) && ({row_reg, col_reg}<18'b001111110010100100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001111110010100100)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001111110010100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b001111110010100110) && ({row_reg, col_reg}<18'b001111110010101000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b001111110010101000) && ({row_reg, col_reg}<18'b001111110010101101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b001111110010101101) && ({row_reg, col_reg}<18'b001111110010101111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b001111110010101111)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001111110010110000)) color_data = 12'b100110111010;
		if(({row_reg, col_reg}==18'b001111110010110001)) color_data = 12'b100110111011;
		if(({row_reg, col_reg}==18'b001111110010110010)) color_data = 12'b100110111100;
		if(({row_reg, col_reg}==18'b001111110010110011)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}==18'b001111110010110100)) color_data = 12'b010001111011;
		if(({row_reg, col_reg}>=18'b001111110010110101) && ({row_reg, col_reg}<18'b001111110010110111)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b001111110010110111)) color_data = 12'b001101111011;
		if(({row_reg, col_reg}==18'b001111110010111000)) color_data = 12'b011010011100;
		if(({row_reg, col_reg}==18'b001111110010111001)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==18'b001111110010111010)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b001111110010111011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001111110010111100)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}>=18'b001111110010111101) && ({row_reg, col_reg}<18'b001111110011000000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001111110011000000) && ({row_reg, col_reg}<18'b001111110011000010)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001111110011000010)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b001111110011000011) && ({row_reg, col_reg}<18'b001111110011001011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001111110011001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001111110011001100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b001111110011001101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001111110011001110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b001111110011001111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001111110011010000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b001111110011010001)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b001111110011010010) && ({row_reg, col_reg}<18'b001111110011010100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b001111110011010100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b001111110011010101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001111110011010110) && ({row_reg, col_reg}<18'b001111110011011001)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b001111110011011001) && ({row_reg, col_reg}<18'b001111110011011101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001111110011011101) && ({row_reg, col_reg}<18'b001111110011100011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001111110011100011)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001111110011100100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001111110011100101)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001111110011100110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001111110011100111) && ({row_reg, col_reg}<18'b001111110011101001)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==18'b001111110011101001)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}>=18'b001111110011101010) && ({row_reg, col_reg}<18'b001111110011101101)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}>=18'b001111110011101101) && ({row_reg, col_reg}<18'b001111110011110000)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}>=18'b001111110011110000) && ({row_reg, col_reg}<18'b001111110011110011)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b001111110011110011) && ({row_reg, col_reg}<18'b001111110011110101)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b001111110011110101) && ({row_reg, col_reg}<18'b001111111000101100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b001111111000101100) && ({row_reg, col_reg}<18'b001111111000110000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b001111111000110000) && ({row_reg, col_reg}<18'b001111111000110010)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}==18'b001111111000110010)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b001111111000110011)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}==18'b001111111000110100)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}>=18'b001111111000110101) && ({row_reg, col_reg}<18'b001111111000110111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001111111000110111) && ({row_reg, col_reg}<18'b001111111000111001)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==18'b001111111000111001)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b001111111000111010) && ({row_reg, col_reg}<18'b001111111000111100)) color_data = 12'b101010111010;
		if(({row_reg, col_reg}==18'b001111111000111100)) color_data = 12'b100111001011;
		if(({row_reg, col_reg}==18'b001111111000111101)) color_data = 12'b101011101101;
		if(({row_reg, col_reg}==18'b001111111000111110)) color_data = 12'b101111101110;
		if(({row_reg, col_reg}==18'b001111111000111111)) color_data = 12'b101111111111;
		if(({row_reg, col_reg}==18'b001111111001000000)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b001111111001000001)) color_data = 12'b010110111101;
		if(({row_reg, col_reg}==18'b001111111001000010)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b001111111001000011)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}>=18'b001111111001000100) && ({row_reg, col_reg}<18'b001111111001001001)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b001111111001001001)) color_data = 12'b001101111011;
		if(({row_reg, col_reg}==18'b001111111001001010)) color_data = 12'b010001111001;
		if(({row_reg, col_reg}==18'b001111111001001011)) color_data = 12'b100110111011;
		if(({row_reg, col_reg}==18'b001111111001001100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001111111001001101)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001111111001001110)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==18'b001111111001001111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b001111111001010000) && ({row_reg, col_reg}<18'b001111111001101000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001111111001101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001111111001101001)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b001111111001101010) && ({row_reg, col_reg}<18'b001111111001101100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001111111001101100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b001111111001101101) && ({row_reg, col_reg}<18'b001111111001110000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001111111001110000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=18'b001111111001110001) && ({row_reg, col_reg}<18'b001111111001110100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001111111001110100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==18'b001111111001110101)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b001111111001110110) && ({row_reg, col_reg}<18'b001111111001111010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001111111001111010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b001111111001111011) && ({row_reg, col_reg}<18'b001111111010000000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001111111010000000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001111111010000001)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b001111111010000010) && ({row_reg, col_reg}<18'b001111111010000100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001111111010000100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001111111010000101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001111111010000110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b001111111010000111) && ({row_reg, col_reg}<18'b001111111010001001)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001111111010001001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001111111010001010) && ({row_reg, col_reg}<18'b001111111010001101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001111111010001101)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b001111111010001110) && ({row_reg, col_reg}<18'b001111111010010010)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001111111010010010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001111111010010011) && ({row_reg, col_reg}<18'b001111111010011011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001111111010011011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001111111010011100) && ({row_reg, col_reg}<18'b001111111010011111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001111111010011111) && ({row_reg, col_reg}<18'b001111111010100001)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b001111111010100001) && ({row_reg, col_reg}<18'b001111111010100011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001111111010100011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b001111111010100100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001111111010100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b001111111010100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001111111010100111)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==18'b001111111010101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001111111010101001) && ({row_reg, col_reg}<18'b001111111010101101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001111111010101101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b001111111010101110)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}==18'b001111111010101111)) color_data = 12'b100110101001;
		if(({row_reg, col_reg}==18'b001111111010110000)) color_data = 12'b100010111001;
		if(({row_reg, col_reg}==18'b001111111010110001)) color_data = 12'b100010111010;
		if(({row_reg, col_reg}==18'b001111111010110010)) color_data = 12'b100110111100;
		if(({row_reg, col_reg}==18'b001111111010110011)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}==18'b001111111010110100)) color_data = 12'b010001111011;
		if(({row_reg, col_reg}>=18'b001111111010110101) && ({row_reg, col_reg}<18'b001111111010110111)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b001111111010110111)) color_data = 12'b001101111011;
		if(({row_reg, col_reg}==18'b001111111010111000)) color_data = 12'b011010011100;
		if(({row_reg, col_reg}==18'b001111111010111001)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==18'b001111111010111010)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}>=18'b001111111010111011) && ({row_reg, col_reg}<18'b001111111010111101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b001111111010111101) && ({row_reg, col_reg}<18'b001111111010111111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001111111010111111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b001111111011000000) && ({row_reg, col_reg}<18'b001111111011000010)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001111111011000010)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b001111111011000011) && ({row_reg, col_reg}<18'b001111111011001001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001111111011001001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001111111011001010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b001111111011001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b001111111011001100) && ({row_reg, col_reg}<18'b001111111011001110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001111111011001110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b001111111011001111) && ({row_reg, col_reg}<18'b001111111011010001)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001111111011010001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001111111011010010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b001111111011010011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b001111111011010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b001111111011010101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b001111111011010110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001111111011010111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001111111011011000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b001111111011011001) && ({row_reg, col_reg}<18'b001111111011011101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001111111011011101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001111111011011110)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b001111111011011111)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==18'b001111111011100000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b001111111011100001)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b001111111011100010)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b001111111011100011) && ({row_reg, col_reg}<18'b001111111011101001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b001111111011101001) && ({row_reg, col_reg}<18'b001111111011101011)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}>=18'b001111111011101011) && ({row_reg, col_reg}<18'b001111111011101101)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}>=18'b001111111011101101) && ({row_reg, col_reg}<18'b001111111011101111)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}==18'b001111111011101111)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}>=18'b001111111011110000) && ({row_reg, col_reg}<18'b001111111011110011)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b001111111011110011) && ({row_reg, col_reg}<18'b001111111011110101)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b001111111011110101) && ({row_reg, col_reg}<18'b010000000000011001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010000000000011001) && ({row_reg, col_reg}<18'b010000000000011011)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010000000000011011) && ({row_reg, col_reg}<18'b010000000000100000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010000000000100000)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}>=18'b010000000000100001) && ({row_reg, col_reg}<18'b010000000000101001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010000000000101001) && ({row_reg, col_reg}<18'b010000000000101101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b010000000000101101)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b010000000000101110) && ({row_reg, col_reg}<18'b010000000000110000)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}==18'b010000000000110000)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}>=18'b010000000000110001) && ({row_reg, col_reg}<18'b010000000000110011)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}>=18'b010000000000110011) && ({row_reg, col_reg}<18'b010000000000110101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000000000110101)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010000000000110110)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}>=18'b010000000000110111) && ({row_reg, col_reg}<18'b010000000000111001)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010000000000111001)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==18'b010000000000111010)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010000000000111011)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}>=18'b010000000000111100) && ({row_reg, col_reg}<18'b010000000000111110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000000000111110)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b010000000000111111)) color_data = 12'b100110111011;
		if(({row_reg, col_reg}==18'b010000000001000000)) color_data = 12'b011111001011;
		if(({row_reg, col_reg}==18'b010000000001000001)) color_data = 12'b100011011101;
		if(({row_reg, col_reg}==18'b010000000001000010)) color_data = 12'b100011011110;
		if(({row_reg, col_reg}==18'b010000000001000011)) color_data = 12'b011111011110;
		if(({row_reg, col_reg}>=18'b010000000001000100) && ({row_reg, col_reg}<18'b010000000001001001)) color_data = 12'b011011011110;
		if(({row_reg, col_reg}==18'b010000000001001001)) color_data = 12'b100011011110;
		if(({row_reg, col_reg}==18'b010000000001001010)) color_data = 12'b100111001101;
		if(({row_reg, col_reg}==18'b010000000001001011)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b010000000001001100)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b010000000001001101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000000001001110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000000001001111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010000000001010000)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010000000001010001) && ({row_reg, col_reg}<18'b010000000001010110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010000000001010110)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==18'b010000000001010111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010000000001011000)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}>=18'b010000000001011001) && ({row_reg, col_reg}<18'b010000000001100111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010000000001100111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010000000001101000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010000000001101001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010000000001101010) && ({row_reg, col_reg}<18'b010000000001101100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010000000001101100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010000000001101101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000000001101110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000000001101111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000000001110000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010000000001110001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010000000001110010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010000000001110011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010000000001110100)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010000000001110101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010000000001110110)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010000000001110111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b010000000001111000) && ({row_reg, col_reg}<18'b010000000001111100)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010000000001111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010000000001111101) && ({row_reg, col_reg}<18'b010000000001111111)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010000000001111111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010000000010000000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010000000010000001) && ({row_reg, col_reg}<18'b010000000010000100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000000010000100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010000000010000101) && ({row_reg, col_reg}<18'b010000000010001000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010000000010001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010000000010001001)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b010000000010001010) && ({row_reg, col_reg}<18'b010000000010001100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010000000010001100)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010000000010001101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010000000010001110) && ({row_reg, col_reg}<18'b010000000010011100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000000010011100)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b010000000010011101) && ({row_reg, col_reg}<18'b010000000010011111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010000000010011111)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010000000010100000)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}>=18'b010000000010100001) && ({row_reg, col_reg}<18'b010000000010100011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010000000010100011) && ({row_reg, col_reg}<18'b010000000010100101)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010000000010100101)) color_data = 12'b100110001001;
		if(({row_reg, col_reg}>=18'b010000000010100110) && ({row_reg, col_reg}<18'b010000000010101000)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010000000010101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010000000010101001) && ({row_reg, col_reg}<18'b010000000010101011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010000000010101011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010000000010101100)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}==18'b010000000010101101)) color_data = 12'b100110101001;
		if(({row_reg, col_reg}==18'b010000000010101110)) color_data = 12'b100010101001;
		if(({row_reg, col_reg}==18'b010000000010101111)) color_data = 12'b101011011100;
		if(({row_reg, col_reg}==18'b010000000010110000)) color_data = 12'b100111101100;
		if(({row_reg, col_reg}==18'b010000000010110001)) color_data = 12'b101011101101;
		if(({row_reg, col_reg}==18'b010000000010110010)) color_data = 12'b101011101111;
		if(({row_reg, col_reg}==18'b010000000010110011)) color_data = 12'b011111001110;
		if(({row_reg, col_reg}==18'b010000000010110100)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b010000000010110101)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010000000010110110)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010000000010110111)) color_data = 12'b010001111100;
		if(({row_reg, col_reg}==18'b010000000010111000)) color_data = 12'b011110001100;
		if(({row_reg, col_reg}==18'b010000000010111001)) color_data = 12'b101010101100;
		if(({row_reg, col_reg}==18'b010000000010111010)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==18'b010000000010111011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000000010111100)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==18'b010000000010111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010000000010111110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010000000010111111)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010000000011000000)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010000000011000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010000000011000010) && ({row_reg, col_reg}<18'b010000000011000101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010000000011000101) && ({row_reg, col_reg}<18'b010000000011001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010000000011001000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010000000011001001) && ({row_reg, col_reg}<18'b010000000011001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010000000011001011)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010000000011001100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010000000011001101) && ({row_reg, col_reg}<18'b010000000011001111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010000000011001111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010000000011010000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010000000011010001) && ({row_reg, col_reg}<18'b010000000011010100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010000000011010100)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}>=18'b010000000011010101) && ({row_reg, col_reg}<18'b010000000011011001)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b010000000011011001) && ({row_reg, col_reg}<18'b010000000011011011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010000000011011011) && ({row_reg, col_reg}<18'b010000000011011110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000000011011110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010000000011011111)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b010000000011100000) && ({row_reg, col_reg}<18'b010000000011100010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010000000011100010)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=18'b010000000011100011) && ({row_reg, col_reg}<18'b010000000011101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010000000011101000) && ({row_reg, col_reg}<18'b010000000011101011)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b010000000011101011) && ({row_reg, col_reg}<18'b010000000011101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010000000011101110)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}==18'b010000000011101111)) color_data = 12'b011110001001;
		if(({row_reg, col_reg}==18'b010000000011110000)) color_data = 12'b011010001010;
		if(({row_reg, col_reg}==18'b010000000011110001)) color_data = 12'b011110011011;
		if(({row_reg, col_reg}==18'b010000000011110010)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b010000000011110011) && ({row_reg, col_reg}<18'b010000000011110101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b010000000011110101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010000000011110110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010000000011110111) && ({row_reg, col_reg}<18'b010000000011111111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010000000011111111)) color_data = 12'b011010101111;

		if(({row_reg, col_reg}>=18'b010000000100000000) && ({row_reg, col_reg}<18'b010000001000011001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010000001000011001)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010000001000011010) && ({row_reg, col_reg}<18'b010000001000101000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010000001000101000) && ({row_reg, col_reg}<18'b010000001000101100)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b010000001000101100)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b010000001000101101) && ({row_reg, col_reg}<18'b010000001000101111)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}==18'b010000001000101111)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}>=18'b010000001000110000) && ({row_reg, col_reg}<18'b010000001000110011)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b010000001000110011)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b010000001000110100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000001000110101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000001000110110)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}>=18'b010000001000110111) && ({row_reg, col_reg}<18'b010000001000111011)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010000001000111011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b010000001000111100) && ({row_reg, col_reg}<18'b010000001000111110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000001000111110)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==18'b010000001000111111)) color_data = 12'b100010011010;
		if(({row_reg, col_reg}==18'b010000001001000000)) color_data = 12'b011110101010;
		if(({row_reg, col_reg}==18'b010000001001000001)) color_data = 12'b100111011101;
		if(({row_reg, col_reg}>=18'b010000001001000010) && ({row_reg, col_reg}<18'b010000001001000100)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}>=18'b010000001001000100) && ({row_reg, col_reg}<18'b010000001001001001)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010000001001001001)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}==18'b010000001001001010)) color_data = 12'b101111101111;
		if(({row_reg, col_reg}==18'b010000001001001011)) color_data = 12'b100110111011;
		if(({row_reg, col_reg}==18'b010000001001001100)) color_data = 12'b101010111011;
		if(({row_reg, col_reg}==18'b010000001001001101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000001001001110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000001001001111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010000001001010000)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010000001001010001) && ({row_reg, col_reg}<18'b010000001001100111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010000001001100111)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010000001001101000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000001001101001)) color_data = 12'b110010111011;
		if(({row_reg, col_reg}>=18'b010000001001101010) && ({row_reg, col_reg}<18'b010000001001101100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==18'b010000001001101100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000001001101101)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}>=18'b010000001001101110) && ({row_reg, col_reg}<18'b010000001001110000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000001001110000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000001001110001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010000001001110010) && ({row_reg, col_reg}<18'b010000001001110100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010000001001110100)) color_data = 12'b011001010101;
		if(({row_reg, col_reg}==18'b010000001001110101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010000001001110110)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010000001001110111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000001001111000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010000001001111001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000001001111010)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010000001001111011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010000001001111100) && ({row_reg, col_reg}<18'b010000001001111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010000001001111110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010000001001111111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b010000001010000000) && ({row_reg, col_reg}<18'b010000001010000011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000001010000011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000001010000100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010000001010000101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010000001010000110) && ({row_reg, col_reg}<18'b010000001010001000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010000001010001000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010000001010001001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010000001010001010) && ({row_reg, col_reg}<18'b010000001010001100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000001010001100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010000001010001101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000001010001110)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}>=18'b010000001010001111) && ({row_reg, col_reg}<18'b010000001010011100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000001010011100)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b010000001010011101) && ({row_reg, col_reg}<18'b010000001010100000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010000001010100000)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==18'b010000001010100001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010000001010100010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010000001010100011) && ({row_reg, col_reg}<18'b010000001010100101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010000001010100101)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010000001010100110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010000001010100111) && ({row_reg, col_reg}<18'b010000001010101010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000001010101010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000001010101011)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==18'b010000001010101100)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b010000001010101101)) color_data = 12'b101010111010;
		if(({row_reg, col_reg}==18'b010000001010101110)) color_data = 12'b100110111010;
		if(({row_reg, col_reg}==18'b010000001010101111)) color_data = 12'b101111101101;
		if(({row_reg, col_reg}==18'b010000001010110000)) color_data = 12'b101011111101;
		if(({row_reg, col_reg}==18'b010000001010110001)) color_data = 12'b101011111110;
		if(({row_reg, col_reg}==18'b010000001010110010)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}==18'b010000001010110011)) color_data = 12'b100011011111;
		if(({row_reg, col_reg}==18'b010000001010110100)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b010000001010110101)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010000001010110110)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010000001010110111)) color_data = 12'b010001111011;
		if(({row_reg, col_reg}==18'b010000001010111000)) color_data = 12'b011110011100;
		if(({row_reg, col_reg}==18'b010000001010111001)) color_data = 12'b101010101100;
		if(({row_reg, col_reg}==18'b010000001010111010)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b010000001010111011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000001010111100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000001010111101)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010000001010111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010000001010111111) && ({row_reg, col_reg}<18'b010000001011000001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010000001011000001)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b010000001011000010) && ({row_reg, col_reg}<18'b010000001011000110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010000001011000110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010000001011000111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010000001011001000) && ({row_reg, col_reg}<18'b010000001011001110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010000001011001110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010000001011001111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010000001011010000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010000001011010001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=18'b010000001011010010) && ({row_reg, col_reg}<18'b010000001011010100)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==18'b010000001011010100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000001011010101)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=18'b010000001011010110) && ({row_reg, col_reg}<18'b010000001011011001)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000001011011001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010000001011011010) && ({row_reg, col_reg}<18'b010000001011011110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000001011011110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010000001011011111)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b010000001011100000) && ({row_reg, col_reg}<18'b010000001011100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010000001011100100) && ({row_reg, col_reg}<18'b010000001011100110)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}>=18'b010000001011100110) && ({row_reg, col_reg}<18'b010000001011101011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010000001011101011) && ({row_reg, col_reg}<18'b010000001011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010000001011101101) && ({row_reg, col_reg}<18'b010000001011110000)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==18'b010000001011110000)) color_data = 12'b011010001010;
		if(({row_reg, col_reg}==18'b010000001011110001)) color_data = 12'b011010011011;
		if(({row_reg, col_reg}==18'b010000001011110010)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b010000001011110011) && ({row_reg, col_reg}<18'b010000001011110101)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b010000001011110101) && ({row_reg, col_reg}<18'b010000010000100000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010000010000100000) && ({row_reg, col_reg}<18'b010000010000100100)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010000010000100100) && ({row_reg, col_reg}<18'b010000010000100111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010000010000100111)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010000010000101000) && ({row_reg, col_reg}<18'b010000010000101011)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b010000010000101011) && ({row_reg, col_reg}<18'b010000010000101101)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}>=18'b010000010000101101) && ({row_reg, col_reg}<18'b010000010000110000)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b010000010000110000)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b010000010000110001)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==18'b010000010000110010)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}==18'b010000010000110011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010000010000110100) && ({row_reg, col_reg}<18'b010000010000111100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000010000111100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000010000111101)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}==18'b010000010000111110)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==18'b010000010000111111)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}==18'b010000010001000000)) color_data = 12'b100010101010;
		if(({row_reg, col_reg}==18'b010000010001000001)) color_data = 12'b101011011100;
		if(({row_reg, col_reg}==18'b010000010001000010)) color_data = 12'b101111101110;
		if(({row_reg, col_reg}==18'b010000010001000011)) color_data = 12'b101011101110;
		if(({row_reg, col_reg}==18'b010000010001000100)) color_data = 12'b100111111110;
		if(({row_reg, col_reg}>=18'b010000010001000101) && ({row_reg, col_reg}<18'b010000010001001000)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010000010001001000)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010000010001001001)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b010000010001001010)) color_data = 12'b101011101110;
		if(({row_reg, col_reg}==18'b010000010001001011)) color_data = 12'b100010111011;
		if(({row_reg, col_reg}==18'b010000010001001100)) color_data = 12'b101010111010;
		if(({row_reg, col_reg}==18'b010000010001001101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000010001001110)) color_data = 12'b101010111010;
		if(({row_reg, col_reg}==18'b010000010001001111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010000010001010000)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}>=18'b010000010001010001) && ({row_reg, col_reg}<18'b010000010001010011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010000010001010011) && ({row_reg, col_reg}<18'b010000010001010101)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010000010001010101) && ({row_reg, col_reg}<18'b010000010001011100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010000010001011100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010000010001011101) && ({row_reg, col_reg}<18'b010000010001100111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010000010001100111)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b010000010001101000) && ({row_reg, col_reg}<18'b010000010001101010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000010001101010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000010001101011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000010001101100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010000010001101101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000010001101110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000010001101111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==18'b010000010001110000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000010001110001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010000010001110010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010000010001110011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010000010001110100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010000010001110101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010000010001110110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010000010001110111)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010000010001111000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010000010001111001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000010001111010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b010000010001111011) && ({row_reg, col_reg}<18'b010000010001111111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010000010001111111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b010000010010000000) && ({row_reg, col_reg}<18'b010000010010000100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000010010000100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010000010010000101) && ({row_reg, col_reg}<18'b010000010010001000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010000010010001000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010000010010001001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b010000010010001010) && ({row_reg, col_reg}<18'b010000010010001110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010000010010001110) && ({row_reg, col_reg}<18'b010000010010011011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b010000010010011011) && ({row_reg, col_reg}<18'b010000010010011101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010000010010011101) && ({row_reg, col_reg}<18'b010000010010011111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010000010010011111)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010000010010100000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010000010010100001)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010000010010100010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010000010010100011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010000010010100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010000010010100101)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b010000010010100110) && ({row_reg, col_reg}<18'b010000010010101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000010010101000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010000010010101001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010000010010101010)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==18'b010000010010101011)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==18'b010000010010101100)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b010000010010101101)) color_data = 12'b101010111011;
		if(({row_reg, col_reg}==18'b010000010010101110)) color_data = 12'b100110111011;
		if(({row_reg, col_reg}==18'b010000010010101111)) color_data = 12'b101111101101;
		if(({row_reg, col_reg}==18'b010000010010110000)) color_data = 12'b101011101101;
		if(({row_reg, col_reg}==18'b010000010010110001)) color_data = 12'b100111101110;
		if(({row_reg, col_reg}==18'b010000010010110010)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b010000010010110011)) color_data = 12'b100011011111;
		if(({row_reg, col_reg}==18'b010000010010110100)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}>=18'b010000010010110101) && ({row_reg, col_reg}<18'b010000010010110111)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010000010010110111)) color_data = 12'b010001101011;
		if(({row_reg, col_reg}==18'b010000010010111000)) color_data = 12'b011110001011;
		if(({row_reg, col_reg}==18'b010000010010111001)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b010000010010111010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010000010010111011) && ({row_reg, col_reg}<18'b010000010010111101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000010010111101)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010000010010111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010000010010111111)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}==18'b010000010011000000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010000010011000001)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b010000010011000010) && ({row_reg, col_reg}<18'b010000010011000110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010000010011000110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010000010011000111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010000010011001000) && ({row_reg, col_reg}<18'b010000010011001010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010000010011001010) && ({row_reg, col_reg}<18'b010000010011001100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010000010011001100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010000010011001101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010000010011001110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010000010011001111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010000010011010000)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==18'b010000010011010001)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000010011010010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000010011010011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b010000010011010100) && ({row_reg, col_reg}<18'b010000010011010111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000010011010111)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b010000010011011000) && ({row_reg, col_reg}<18'b010000010011011110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000010011011110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010000010011011111)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b010000010011100000) && ({row_reg, col_reg}<18'b010000010011100010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010000010011100010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010000010011100011) && ({row_reg, col_reg}<18'b010000010011100101)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}>=18'b010000010011100101) && ({row_reg, col_reg}<18'b010000010011101011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010000010011101011) && ({row_reg, col_reg}<18'b010000010011101101)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010000010011101101)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==18'b010000010011101110)) color_data = 12'b011110001000;
		if(({row_reg, col_reg}==18'b010000010011101111)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==18'b010000010011110000)) color_data = 12'b010110001001;
		if(({row_reg, col_reg}==18'b010000010011110001)) color_data = 12'b011010001011;
		if(({row_reg, col_reg}==18'b010000010011110010)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}>=18'b010000010011110011) && ({row_reg, col_reg}<18'b010000010011110101)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b010000010011110101) && ({row_reg, col_reg}<18'b010000011000100000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010000011000100000) && ({row_reg, col_reg}<18'b010000011000100011)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b010000011000100011)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}>=18'b010000011000100100) && ({row_reg, col_reg}<18'b010000011000100111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010000011000100111)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010000011000101000) && ({row_reg, col_reg}<18'b010000011000101010)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b010000011000101010)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}>=18'b010000011000101011) && ({row_reg, col_reg}<18'b010000011000101110)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}>=18'b010000011000101110) && ({row_reg, col_reg}<18'b010000011000110000)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}==18'b010000011000110000)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}>=18'b010000011000110001) && ({row_reg, col_reg}<18'b010000011000110011)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}==18'b010000011000110011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010000011000110100) && ({row_reg, col_reg}<18'b010000011000111100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000011000111100)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}>=18'b010000011000111101) && ({row_reg, col_reg}<18'b010000011000111111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010000011000111111) && ({row_reg, col_reg}<18'b010000011001000001)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==18'b010000011001000001)) color_data = 12'b101111001100;
		if(({row_reg, col_reg}==18'b010000011001000010)) color_data = 12'b110011101110;
		if(({row_reg, col_reg}==18'b010000011001000011)) color_data = 12'b101111101110;
		if(({row_reg, col_reg}==18'b010000011001000100)) color_data = 12'b101011111110;
		if(({row_reg, col_reg}==18'b010000011001000101)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}>=18'b010000011001000110) && ({row_reg, col_reg}<18'b010000011001001010)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010000011001001010)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}==18'b010000011001001011)) color_data = 12'b100011001100;
		if(({row_reg, col_reg}==18'b010000011001001100)) color_data = 12'b100110111011;
		if(({row_reg, col_reg}>=18'b010000011001001101) && ({row_reg, col_reg}<18'b010000011001001111)) color_data = 12'b101010111011;
		if(({row_reg, col_reg}==18'b010000011001001111)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}>=18'b010000011001010000) && ({row_reg, col_reg}<18'b010000011001010010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010000011001010010) && ({row_reg, col_reg}<18'b010000011001010101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010000011001010101)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010000011001010110) && ({row_reg, col_reg}<18'b010000011001011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010000011001011000) && ({row_reg, col_reg}<18'b010000011001011010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010000011001011010) && ({row_reg, col_reg}<18'b010000011001011100)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==18'b010000011001011100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010000011001011101)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010000011001011110) && ({row_reg, col_reg}<18'b010000011001100000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010000011001100000) && ({row_reg, col_reg}<18'b010000011001100010)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010000011001100010) && ({row_reg, col_reg}<18'b010000011001100100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010000011001100100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010000011001100101) && ({row_reg, col_reg}<18'b010000011001100111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010000011001100111)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b010000011001101000) && ({row_reg, col_reg}<18'b010000011001101111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000011001101111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==18'b010000011001110000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000011001110001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010000011001110010) && ({row_reg, col_reg}<18'b010000011001110101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010000011001110101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010000011001110110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010000011001110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010000011001111000) && ({row_reg, col_reg}<18'b010000011001111011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010000011001111011) && ({row_reg, col_reg}<18'b010000011001111111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010000011001111111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010000011010000000) && ({row_reg, col_reg}<18'b010000011010000011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000011010000011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000011010000100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010000011010000101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010000011010000110) && ({row_reg, col_reg}<18'b010000011010001000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010000011010001000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010000011010001001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b010000011010001010) && ({row_reg, col_reg}<18'b010000011010001101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010000011010001101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010000011010001110) && ({row_reg, col_reg}<18'b010000011010011011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000011010011011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000011010011100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000011010011101)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010000011010011110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010000011010011111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000011010100000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010000011010100001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010000011010100010) && ({row_reg, col_reg}<18'b010000011010100101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010000011010100101)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010000011010100110)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010000011010100111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010000011010101000) && ({row_reg, col_reg}<18'b010000011010101010)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010000011010101010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000011010101011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000011010101100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000011010101101)) color_data = 12'b101010111011;
		if(({row_reg, col_reg}==18'b010000011010101110)) color_data = 12'b100110111011;
		if(({row_reg, col_reg}==18'b010000011010101111)) color_data = 12'b101011101110;
		if(({row_reg, col_reg}==18'b010000011010110000)) color_data = 12'b100111101110;
		if(({row_reg, col_reg}>=18'b010000011010110001) && ({row_reg, col_reg}<18'b010000011010110011)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}==18'b010000011010110011)) color_data = 12'b100011011111;
		if(({row_reg, col_reg}>=18'b010000011010110100) && ({row_reg, col_reg}<18'b010000011010110110)) color_data = 12'b001101111011;
		if(({row_reg, col_reg}==18'b010000011010110110)) color_data = 12'b010001101011;
		if(({row_reg, col_reg}==18'b010000011010110111)) color_data = 12'b010001101001;
		if(({row_reg, col_reg}==18'b010000011010111000)) color_data = 12'b011110001011;
		if(({row_reg, col_reg}==18'b010000011010111001)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b010000011010111010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010000011010111011) && ({row_reg, col_reg}<18'b010000011010111101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000011010111101)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010000011010111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010000011010111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010000011011000000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010000011011000001)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b010000011011000010) && ({row_reg, col_reg}<18'b010000011011000110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010000011011000110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010000011011000111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010000011011001000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010000011011001001) && ({row_reg, col_reg}<18'b010000011011001011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010000011011001011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010000011011001100) && ({row_reg, col_reg}<18'b010000011011001110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010000011011001110) && ({row_reg, col_reg}<18'b010000011011010000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010000011011010000)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010000011011010001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==18'b010000011011010010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010000011011010011) && ({row_reg, col_reg}<18'b010000011011010110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000011011010110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000011011010111)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}>=18'b010000011011011000) && ({row_reg, col_reg}<18'b010000011011011100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000011011011100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==18'b010000011011011101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000011011011110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010000011011011111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010000011011100000) && ({row_reg, col_reg}<18'b010000011011100010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010000011011100010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010000011011100011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010000011011100100)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}>=18'b010000011011100101) && ({row_reg, col_reg}<18'b010000011011101101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010000011011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010000011011101110) && ({row_reg, col_reg}<18'b010000011011110000)) color_data = 12'b011110001000;
		if(({row_reg, col_reg}==18'b010000011011110000)) color_data = 12'b011010001001;
		if(({row_reg, col_reg}==18'b010000011011110001)) color_data = 12'b011010001011;
		if(({row_reg, col_reg}==18'b010000011011110010)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}==18'b010000011011110011)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b010000011011110100)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010000011011110101) && ({row_reg, col_reg}<18'b010000011011111101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010000011011111101) && ({row_reg, col_reg}<18'b010000011100000000)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b010000011100000000) && ({row_reg, col_reg}<18'b010000100000100000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010000100000100000) && ({row_reg, col_reg}<18'b010000100000100010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010000100000100010) && ({row_reg, col_reg}<18'b010000100000100100)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}>=18'b010000100000100100) && ({row_reg, col_reg}<18'b010000100000100111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010000100000100111)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}>=18'b010000100000101000) && ({row_reg, col_reg}<18'b010000100000101010)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b010000100000101010) && ({row_reg, col_reg}<18'b010000100000101100)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b010000100000101100)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}>=18'b010000100000101101) && ({row_reg, col_reg}<18'b010000100000110000)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}>=18'b010000100000110000) && ({row_reg, col_reg}<18'b010000100000110011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010000100000110011) && ({row_reg, col_reg}<18'b010000100000110111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000100000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000100000111000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010000100000111001)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b010000100000111010) && ({row_reg, col_reg}<18'b010000100000111101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000100000111101)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==18'b010000100000111110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b010000100000111111) && ({row_reg, col_reg}<18'b010000100001000001)) color_data = 12'b100010011000;
		if(({row_reg, col_reg}==18'b010000100001000001)) color_data = 12'b101010111010;
		if(({row_reg, col_reg}>=18'b010000100001000010) && ({row_reg, col_reg}<18'b010000100001000100)) color_data = 12'b101111011100;
		if(({row_reg, col_reg}==18'b010000100001000100)) color_data = 12'b101011011101;
		if(({row_reg, col_reg}==18'b010000100001000101)) color_data = 12'b101011101110;
		if(({row_reg, col_reg}==18'b010000100001000110)) color_data = 12'b100011011110;
		if(({row_reg, col_reg}==18'b010000100001000111)) color_data = 12'b011111011110;
		if(({row_reg, col_reg}>=18'b010000100001001000) && ({row_reg, col_reg}<18'b010000100001001010)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}==18'b010000100001001010)) color_data = 12'b100011011111;
		if(({row_reg, col_reg}==18'b010000100001001011)) color_data = 12'b011110111101;
		if(({row_reg, col_reg}==18'b010000100001001100)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}==18'b010000100001001101)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}>=18'b010000100001001110) && ({row_reg, col_reg}<18'b010000100001010000)) color_data = 12'b100010011011;
		if(({row_reg, col_reg}>=18'b010000100001010000) && ({row_reg, col_reg}<18'b010000100001010011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010000100001010011)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010000100001010100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010000100001010101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010000100001010110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010000100001010111) && ({row_reg, col_reg}<18'b010000100001011001)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010000100001011001) && ({row_reg, col_reg}<18'b010000100001011100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010000100001011100) && ({row_reg, col_reg}<18'b010000100001011110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010000100001011110) && ({row_reg, col_reg}<18'b010000100001100000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010000100001100000) && ({row_reg, col_reg}<18'b010000100001100011)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==18'b010000100001100011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010000100001100100) && ({row_reg, col_reg}<18'b010000100001100110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010000100001100110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010000100001100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010000100001101000) && ({row_reg, col_reg}<18'b010000100001101100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b010000100001101100) && ({row_reg, col_reg}<18'b010000100001101110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000100001101110)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==18'b010000100001101111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000100001110000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010000100001110001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010000100001110010) && ({row_reg, col_reg}<18'b010000100001110101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010000100001110101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010000100001110110)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b010000100001110111) && ({row_reg, col_reg}<18'b010000100001111001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b010000100001111001) && ({row_reg, col_reg}<18'b010000100001111011)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b010000100001111011) && ({row_reg, col_reg}<18'b010000100001111111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010000100001111111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010000100010000000) && ({row_reg, col_reg}<18'b010000100010000100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000100010000100)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b010000100010000101) && ({row_reg, col_reg}<18'b010000100010001000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010000100010001000)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010000100010001001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010000100010001010) && ({row_reg, col_reg}<18'b010000100010001101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000100010001101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000100010001110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010000100010001111) && ({row_reg, col_reg}<18'b010000100010011000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000100010011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000100010011001)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000100010011010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010000100010011011) && ({row_reg, col_reg}<18'b010000100010011101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010000100010011101)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010000100010011110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010000100010011111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010000100010100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010000100010100001) && ({row_reg, col_reg}<18'b010000100010100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010000100010100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010000100010100110)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010000100010100111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010000100010101000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010000100010101001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010000100010101010)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==18'b010000100010101011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000100010101100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000100010101101)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b010000100010101110)) color_data = 12'b100110111100;
		if(({row_reg, col_reg}==18'b010000100010101111)) color_data = 12'b100010111101;
		if(({row_reg, col_reg}==18'b010000100010110000)) color_data = 12'b011111001101;
		if(({row_reg, col_reg}==18'b010000100010110001)) color_data = 12'b011111011110;
		if(({row_reg, col_reg}==18'b010000100010110010)) color_data = 12'b011111001111;
		if(({row_reg, col_reg}==18'b010000100010110011)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==18'b010000100010110100)) color_data = 12'b010010001011;
		if(({row_reg, col_reg}==18'b010000100010110101)) color_data = 12'b010110001100;
		if(({row_reg, col_reg}==18'b010000100010110110)) color_data = 12'b011010001011;
		if(({row_reg, col_reg}==18'b010000100010110111)) color_data = 12'b011001111010;
		if(({row_reg, col_reg}==18'b010000100010111000)) color_data = 12'b100010011011;
		if(({row_reg, col_reg}==18'b010000100010111001)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}>=18'b010000100010111010) && ({row_reg, col_reg}<18'b010000100010111100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000100010111100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000100010111101)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b010000100010111110) && ({row_reg, col_reg}<18'b010000100011000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010000100011000000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010000100011000001)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010000100011000010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010000100011000011) && ({row_reg, col_reg}<18'b010000100011000101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010000100011000101)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010000100011000110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010000100011000111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010000100011001000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010000100011001001) && ({row_reg, col_reg}<18'b010000100011001011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010000100011001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010000100011001100)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010000100011001101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010000100011001110)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010000100011001111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010000100011010000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010000100011010001)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000100011010010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010000100011010011) && ({row_reg, col_reg}<18'b010000100011010110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000100011010110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010000100011010111) && ({row_reg, col_reg}<18'b010000100011011001)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000100011011001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010000100011011010) && ({row_reg, col_reg}<18'b010000100011011101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010000100011011101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010000100011011110)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b010000100011011111) && ({row_reg, col_reg}<18'b010000100011100010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010000100011100010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010000100011100011)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}==18'b010000100011100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010000100011100101)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}==18'b010000100011100110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010000100011100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010000100011101000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010000100011101001) && ({row_reg, col_reg}<18'b010000100011101011)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==18'b010000100011101011)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010000100011101100) && ({row_reg, col_reg}<18'b010000100011101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010000100011101110)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==18'b010000100011101111)) color_data = 12'b011110001000;
		if(({row_reg, col_reg}==18'b010000100011110000)) color_data = 12'b011001111001;
		if(({row_reg, col_reg}==18'b010000100011110001)) color_data = 12'b011010001010;
		if(({row_reg, col_reg}==18'b010000100011110010)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}>=18'b010000100011110011) && ({row_reg, col_reg}<18'b010000100011110101)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b010000100011110101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010000100011110110) && ({row_reg, col_reg}<18'b010000100011111101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010000100011111101) && ({row_reg, col_reg}<18'b010000100100000000)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b010000100100000000) && ({row_reg, col_reg}<18'b010000101000010000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010000101000010000) && ({row_reg, col_reg}<18'b010000101000010010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010000101000010010) && ({row_reg, col_reg}<18'b010000101000100000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010000101000100000)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}==18'b010000101000100001)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010000101000100010) && ({row_reg, col_reg}<18'b010000101000100100)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}==18'b010000101000100100)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b010000101000100101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010000101000100110)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==18'b010000101000100111)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}==18'b010000101000101000)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b010000101000101001)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}==18'b010000101000101010)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b010000101000101011)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}>=18'b010000101000101100) && ({row_reg, col_reg}<18'b010000101000101111)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b010000101000101111)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}>=18'b010000101000110000) && ({row_reg, col_reg}<18'b010000101000110011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010000101000110011) && ({row_reg, col_reg}<18'b010000101000111000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000101000111000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000101000111001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010000101000111010)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010000101000111011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010000101000111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010000101000111101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010000101000111110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010000101000111111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010000101001000000)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==18'b010000101001000001)) color_data = 12'b100010011000;
		if(({row_reg, col_reg}==18'b010000101001000010)) color_data = 12'b101010111010;
		if(({row_reg, col_reg}==18'b010000101001000011)) color_data = 12'b100110111011;
		if(({row_reg, col_reg}==18'b010000101001000100)) color_data = 12'b100110111100;
		if(({row_reg, col_reg}==18'b010000101001000101)) color_data = 12'b100010111100;
		if(({row_reg, col_reg}==18'b010000101001000110)) color_data = 12'b010110011011;
		if(({row_reg, col_reg}==18'b010000101001000111)) color_data = 12'b001110001011;
		if(({row_reg, col_reg}==18'b010000101001001000)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b010000101001001001)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b010000101001001010)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b010000101001001011)) color_data = 12'b001101111011;
		if(({row_reg, col_reg}>=18'b010000101001001100) && ({row_reg, col_reg}<18'b010000101001001110)) color_data = 12'b010001111011;
		if(({row_reg, col_reg}==18'b010000101001001110)) color_data = 12'b010101111010;
		if(({row_reg, col_reg}==18'b010000101001001111)) color_data = 12'b011010001011;
		if(({row_reg, col_reg}==18'b010000101001010000)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}>=18'b010000101001010001) && ({row_reg, col_reg}<18'b010000101001010011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000101001010011)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==18'b010000101001010100)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010000101001010101)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010000101001010110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010000101001010111)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010000101001011000) && ({row_reg, col_reg}<18'b010000101001011010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010000101001011010) && ({row_reg, col_reg}<18'b010000101001011100)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}>=18'b010000101001011100) && ({row_reg, col_reg}<18'b010000101001011110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010000101001011110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010000101001011111)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==18'b010000101001100000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010000101001100001) && ({row_reg, col_reg}<18'b010000101001100011)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==18'b010000101001100011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010000101001100100) && ({row_reg, col_reg}<18'b010000101001100110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010000101001100110)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}==18'b010000101001100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010000101001101000) && ({row_reg, col_reg}<18'b010000101001101101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000101001101101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000101001101110)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==18'b010000101001101111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000101001110000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010000101001110001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010000101001110010) && ({row_reg, col_reg}<18'b010000101001110110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010000101001110110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010000101001110111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010000101001111000) && ({row_reg, col_reg}<18'b010000101001111101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010000101001111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010000101001111110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010000101001111111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010000101010000000) && ({row_reg, col_reg}<18'b010000101010000100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000101010000100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010000101010000101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b010000101010000110) && ({row_reg, col_reg}<18'b010000101010001001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010000101010001001) && ({row_reg, col_reg}<18'b010000101010001100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000101010001100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010000101010001101) && ({row_reg, col_reg}<18'b010000101010010111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000101010010111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000101010011000)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010000101010011001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010000101010011010)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010000101010011011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010000101010011100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010000101010011101) && ({row_reg, col_reg}<18'b010000101010011111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010000101010011111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010000101010100000)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}==18'b010000101010100001)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010000101010100010) && ({row_reg, col_reg}<18'b010000101010100100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010000101010100100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010000101010100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010000101010100110) && ({row_reg, col_reg}<18'b010000101010101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000101010101000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010000101010101001)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b010000101010101010) && ({row_reg, col_reg}<18'b010000101010101100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000101010101100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000101010101101)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b010000101010101110)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b010000101010101111)) color_data = 12'b010110001010;
		if(({row_reg, col_reg}==18'b010000101010110000)) color_data = 12'b001110001011;
		if(({row_reg, col_reg}>=18'b010000101010110001) && ({row_reg, col_reg}<18'b010000101010110011)) color_data = 12'b001110001010;
		if(({row_reg, col_reg}==18'b010000101010110011)) color_data = 12'b010010011011;
		if(({row_reg, col_reg}==18'b010000101010110100)) color_data = 12'b011010101100;
		if(({row_reg, col_reg}==18'b010000101010110101)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b010000101010110110)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}==18'b010000101010110111)) color_data = 12'b100010011011;
		if(({row_reg, col_reg}==18'b010000101010111000)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}==18'b010000101010111001)) color_data = 12'b101010111011;
		if(({row_reg, col_reg}>=18'b010000101010111010) && ({row_reg, col_reg}<18'b010000101010111100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000101010111100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000101010111101)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b010000101010111110) && ({row_reg, col_reg}<18'b010000101011000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010000101011000001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010000101011000010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010000101011000011) && ({row_reg, col_reg}<18'b010000101011000110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010000101011000110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010000101011000111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010000101011001000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010000101011001001) && ({row_reg, col_reg}<18'b010000101011001011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010000101011001011)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010000101011001100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000101011001101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010000101011001110) && ({row_reg, col_reg}<18'b010000101011010001)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000101011010001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=18'b010000101011010010) && ({row_reg, col_reg}<18'b010000101011010110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000101011010110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010000101011010111) && ({row_reg, col_reg}<18'b010000101011011001)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000101011011001)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010000101011011010)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b010000101011011011) && ({row_reg, col_reg}<18'b010000101011011101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010000101011011101) && ({row_reg, col_reg}<18'b010000101011100100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010000101011100100)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}==18'b010000101011100101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010000101011100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010000101011100111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010000101011101000) && ({row_reg, col_reg}<18'b010000101011101100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010000101011101100) && ({row_reg, col_reg}<18'b010000101011101111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010000101011101111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010000101011110000)) color_data = 12'b011001111001;
		if(({row_reg, col_reg}==18'b010000101011110001)) color_data = 12'b011010001010;
		if(({row_reg, col_reg}==18'b010000101011110010)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}>=18'b010000101011110011) && ({row_reg, col_reg}<18'b010000101011110101)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b010000101011110101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010000101011110110) && ({row_reg, col_reg}<18'b010000101011111101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010000101011111101) && ({row_reg, col_reg}<18'b010000101100000000)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b010000101100000000) && ({row_reg, col_reg}<18'b010000110000100000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010000110000100000)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}==18'b010000110000100001)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010000110000100010) && ({row_reg, col_reg}<18'b010000110000100100)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}==18'b010000110000100100)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b010000110000100101)) color_data = 12'b011010111111;
		if(({row_reg, col_reg}==18'b010000110000100110)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==18'b010000110000100111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010000110000101000)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b010000110000101001)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}==18'b010000110000101010)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b010000110000101011)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}>=18'b010000110000101100) && ({row_reg, col_reg}<18'b010000110000101110)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}>=18'b010000110000101110) && ({row_reg, col_reg}<18'b010000110000110000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010000110000110000) && ({row_reg, col_reg}<18'b010000110000110100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000110000110100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000110000110101)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==18'b010000110000110110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000110000110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010000110000111000) && ({row_reg, col_reg}<18'b010000110000111011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010000110000111011)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010000110000111100)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010000110000111101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010000110000111110) && ({row_reg, col_reg}<18'b010000110001000000)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010000110001000000)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==18'b010000110001000001)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==18'b010000110001000010)) color_data = 12'b101010111011;
		if(({row_reg, col_reg}==18'b010000110001000011)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b010000110001000100)) color_data = 12'b100110111100;
		if(({row_reg, col_reg}==18'b010000110001000101)) color_data = 12'b100010111101;
		if(({row_reg, col_reg}==18'b010000110001000110)) color_data = 12'b010110001011;
		if(({row_reg, col_reg}==18'b010000110001000111)) color_data = 12'b001101111010;
		if(({row_reg, col_reg}==18'b010000110001001000)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010000110001001001)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b010000110001001010) && ({row_reg, col_reg}<18'b010000110001001100)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010000110001001100)) color_data = 12'b010001111101;
		if(({row_reg, col_reg}==18'b010000110001001101)) color_data = 12'b010001111100;
		if(({row_reg, col_reg}==18'b010000110001001110)) color_data = 12'b010001101011;
		if(({row_reg, col_reg}==18'b010000110001001111)) color_data = 12'b010101111011;
		if(({row_reg, col_reg}==18'b010000110001010000)) color_data = 12'b101010111100;
		if(({row_reg, col_reg}==18'b010000110001010001)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b010000110001010010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000110001010011)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==18'b010000110001010100)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}>=18'b010000110001010101) && ({row_reg, col_reg}<18'b010000110001010111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010000110001010111) && ({row_reg, col_reg}<18'b010000110001011001)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010000110001011001) && ({row_reg, col_reg}<18'b010000110001011100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010000110001011100) && ({row_reg, col_reg}<18'b010000110001011110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010000110001011110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010000110001011111)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010000110001100000) && ({row_reg, col_reg}<18'b010000110001100100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010000110001100100) && ({row_reg, col_reg}<18'b010000110001100110)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}==18'b010000110001100110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010000110001100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010000110001101000) && ({row_reg, col_reg}<18'b010000110001101011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000110001101011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010000110001101100) && ({row_reg, col_reg}<18'b010000110001101110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010000110001101110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010000110001101111)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==18'b010000110001110000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b010000110001110001) && ({row_reg, col_reg}<18'b010000110001110011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010000110001110011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010000110001110100) && ({row_reg, col_reg}<18'b010000110001110110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010000110001110110) && ({row_reg, col_reg}<18'b010000110001111000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010000110001111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010000110001111001) && ({row_reg, col_reg}<18'b010000110001111011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010000110001111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010000110001111100)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b010000110001111101) && ({row_reg, col_reg}<18'b010000110001111111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010000110001111111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010000110010000000) && ({row_reg, col_reg}<18'b010000110010000100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b010000110010000100) && ({row_reg, col_reg}<18'b010000110010001000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000110010001000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010000110010001001) && ({row_reg, col_reg}<18'b010000110010010111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000110010010111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010000110010011000) && ({row_reg, col_reg}<18'b010000110010011100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010000110010011100)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010000110010011101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010000110010011110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010000110010011111)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010000110010100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010000110010100001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010000110010100010) && ({row_reg, col_reg}<18'b010000110010100100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010000110010100100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010000110010100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010000110010100110) && ({row_reg, col_reg}<18'b010000110010101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000110010101000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010000110010101001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010000110010101010)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}>=18'b010000110010101011) && ({row_reg, col_reg}<18'b010000110010101101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000110010101101)) color_data = 12'b101010101100;
		if(({row_reg, col_reg}==18'b010000110010101110)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==18'b010000110010101111)) color_data = 12'b010101111010;
		if(({row_reg, col_reg}==18'b010000110010110000)) color_data = 12'b010001111011;
		if(({row_reg, col_reg}==18'b010000110010110001)) color_data = 12'b001101111011;
		if(({row_reg, col_reg}==18'b010000110010110010)) color_data = 12'b001101111010;
		if(({row_reg, col_reg}==18'b010000110010110011)) color_data = 12'b010010001010;
		if(({row_reg, col_reg}==18'b010000110010110100)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}==18'b010000110010110101)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}>=18'b010000110010110110) && ({row_reg, col_reg}<18'b010000110010111001)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==18'b010000110010111001)) color_data = 12'b101010111011;
		if(({row_reg, col_reg}==18'b010000110010111010)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}>=18'b010000110010111011) && ({row_reg, col_reg}<18'b010000110010111101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000110010111101)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b010000110010111110) && ({row_reg, col_reg}<18'b010000110011000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010000110011000000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010000110011000001)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010000110011000010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010000110011000011) && ({row_reg, col_reg}<18'b010000110011000110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010000110011000110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010000110011000111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010000110011001000) && ({row_reg, col_reg}<18'b010000110011001011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010000110011001011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010000110011001100)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}>=18'b010000110011001101) && ({row_reg, col_reg}<18'b010000110011001111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000110011001111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=18'b010000110011010000) && ({row_reg, col_reg}<18'b010000110011010010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000110011010010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000110011010011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000110011010100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010000110011010101) && ({row_reg, col_reg}<18'b010000110011010111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000110011010111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000110011011000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000110011011001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010000110011011010) && ({row_reg, col_reg}<18'b010000110011100100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010000110011100100) && ({row_reg, col_reg}<18'b010000110011100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010000110011100110) && ({row_reg, col_reg}<18'b010000110011101000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010000110011101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010000110011101001) && ({row_reg, col_reg}<18'b010000110011101011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010000110011101011)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==18'b010000110011101100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010000110011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010000110011101110) && ({row_reg, col_reg}<18'b010000110011110000)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010000110011110000)) color_data = 12'b011001111000;
		if(({row_reg, col_reg}==18'b010000110011110001)) color_data = 12'b011110001010;
		if(({row_reg, col_reg}>=18'b010000110011110010) && ({row_reg, col_reg}<18'b010000110011110100)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b010000110011110100)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b010000110011110101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010000110011110110) && ({row_reg, col_reg}<18'b010000110011111101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010000110011111101) && ({row_reg, col_reg}<18'b010000110100000000)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b010000110100000000) && ({row_reg, col_reg}<18'b010000111000011000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010000111000011000) && ({row_reg, col_reg}<18'b010000111000011010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010000111000011010) && ({row_reg, col_reg}<18'b010000111000100001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010000111000100001)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}==18'b010000111000100010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010000111000100011) && ({row_reg, col_reg}<18'b010000111000100101)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b010000111000100101)) color_data = 12'b011010111111;
		if(({row_reg, col_reg}>=18'b010000111000100110) && ({row_reg, col_reg}<18'b010000111000101000)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==18'b010000111000101000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b010000111000101001)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}==18'b010000111000101010)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}>=18'b010000111000101011) && ({row_reg, col_reg}<18'b010000111000101101)) color_data = 12'b100110011011;
		if(({row_reg, col_reg}==18'b010000111000101101)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}>=18'b010000111000101110) && ({row_reg, col_reg}<18'b010000111000110000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010000111000110000) && ({row_reg, col_reg}<18'b010000111000110011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000111000110011)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}>=18'b010000111000110100) && ({row_reg, col_reg}<18'b010000111000111000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000111000111000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010000111000111001) && ({row_reg, col_reg}<18'b010000111000111011)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010000111000111011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000111000111100)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b010000111000111101) && ({row_reg, col_reg}<18'b010000111000111111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010000111000111111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010000111001000000)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}==18'b010000111001000001)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==18'b010000111001000010)) color_data = 12'b101010111011;
		if(({row_reg, col_reg}==18'b010000111001000011)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b010000111001000100)) color_data = 12'b101010111101;
		if(({row_reg, col_reg}==18'b010000111001000101)) color_data = 12'b100110111110;
		if(({row_reg, col_reg}==18'b010000111001000110)) color_data = 12'b011010001100;
		if(({row_reg, col_reg}==18'b010000111001000111)) color_data = 12'b010001111011;
		if(({row_reg, col_reg}==18'b010000111001001000)) color_data = 12'b010001111100;
		if(({row_reg, col_reg}==18'b010000111001001001)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}>=18'b010000111001001010) && ({row_reg, col_reg}<18'b010000111001001100)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010000111001001100)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010000111001001101)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010000111001001110)) color_data = 12'b001101101011;
		if(({row_reg, col_reg}==18'b010000111001001111)) color_data = 12'b010001111011;
		if(({row_reg, col_reg}==18'b010000111001010000)) color_data = 12'b101010111101;
		if(({row_reg, col_reg}==18'b010000111001010001)) color_data = 12'b101010111100;
		if(({row_reg, col_reg}==18'b010000111001010010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000111001010011)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==18'b010000111001010100)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==18'b010000111001010101)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==18'b010000111001010110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010000111001010111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010000111001011000)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010000111001011001) && ({row_reg, col_reg}<18'b010000111001011101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010000111001011101) && ({row_reg, col_reg}<18'b010000111001100100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010000111001100100) && ({row_reg, col_reg}<18'b010000111001100111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010000111001100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010000111001101000) && ({row_reg, col_reg}<18'b010000111001101101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000111001101101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000111001101110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010000111001101111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000111001110000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010000111001110001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010000111001110010) && ({row_reg, col_reg}<18'b010000111001110110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010000111001110110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010000111001110111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010000111001111000) && ({row_reg, col_reg}<18'b010000111001111111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010000111001111111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010000111010000000) && ({row_reg, col_reg}<18'b010000111010000100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b010000111010000100) && ({row_reg, col_reg}<18'b010000111010000111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010000111010000111) && ({row_reg, col_reg}<18'b010000111010001001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010000111010001001) && ({row_reg, col_reg}<18'b010000111010010111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000111010010111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000111010011000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010000111010011001)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b010000111010011010) && ({row_reg, col_reg}<18'b010000111010011100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010000111010011100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010000111010011101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010000111010011110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010000111010011111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010000111010100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010000111010100001) && ({row_reg, col_reg}<18'b010000111010100101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010000111010100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010000111010100110) && ({row_reg, col_reg}<18'b010000111010101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000111010101000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010000111010101001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010000111010101010)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}>=18'b010000111010101011) && ({row_reg, col_reg}<18'b010000111010101101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000111010101101)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b010000111010101110)) color_data = 12'b100110111101;
		if(({row_reg, col_reg}==18'b010000111010101111)) color_data = 12'b010101111010;
		if(({row_reg, col_reg}>=18'b010000111010110000) && ({row_reg, col_reg}<18'b010000111010110010)) color_data = 12'b010001111011;
		if(({row_reg, col_reg}==18'b010000111010110010)) color_data = 12'b010001111010;
		if(({row_reg, col_reg}==18'b010000111010110011)) color_data = 12'b010101111001;
		if(({row_reg, col_reg}==18'b010000111010110100)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b010000111010110101)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==18'b010000111010110110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010000111010110111)) color_data = 12'b100110101001;
		if(({row_reg, col_reg}==18'b010000111010111000)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==18'b010000111010111001)) color_data = 12'b101010111011;
		if(({row_reg, col_reg}>=18'b010000111010111010) && ({row_reg, col_reg}<18'b010000111010111100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010000111010111100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000111010111101)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010000111010111110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010000111010111111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010000111011000000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010000111011000001)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010000111011000010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010000111011000011) && ({row_reg, col_reg}<18'b010000111011000101)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010000111011000101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010000111011000110) && ({row_reg, col_reg}<18'b010000111011001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010000111011001000) && ({row_reg, col_reg}<18'b010000111011001011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010000111011001011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010000111011001100) && ({row_reg, col_reg}<18'b010000111011001110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000111011001110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010000111011001111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b010000111011010000) && ({row_reg, col_reg}<18'b010000111011010010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010000111011010010) && ({row_reg, col_reg}<18'b010000111011010101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000111011010101)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}>=18'b010000111011010110) && ({row_reg, col_reg}<18'b010000111011011000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010000111011011000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==18'b010000111011011001)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b010000111011011010) && ({row_reg, col_reg}<18'b010000111011100011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010000111011100011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010000111011100100) && ({row_reg, col_reg}<18'b010000111011101000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010000111011101000)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010000111011101001) && ({row_reg, col_reg}<18'b010000111011101011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010000111011101011)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==18'b010000111011101100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010000111011101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010000111011101110)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010000111011101111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010000111011110000)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==18'b010000111011110001)) color_data = 12'b011110001001;
		if(({row_reg, col_reg}==18'b010000111011110010)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}==18'b010000111011110011)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b010000111011110100)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}==18'b010000111011110101)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b010000111011110110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010000111011110111) && ({row_reg, col_reg}<18'b010000111011111101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010000111011111101) && ({row_reg, col_reg}<18'b010000111100000000)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b010000111100000000) && ({row_reg, col_reg}<18'b010001000000010010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010001000000010010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010001000000010011) && ({row_reg, col_reg}<18'b010001000000010111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010001000000010111)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b010001000000011000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010001000000011001) && ({row_reg, col_reg}<18'b010001000000011011)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010001000000011011) && ({row_reg, col_reg}<18'b010001000000100001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010001000000100001)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b010001000000100010)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}>=18'b010001000000100011) && ({row_reg, col_reg}<18'b010001000000100110)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b010001000000100110) && ({row_reg, col_reg}<18'b010001000000101000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010001000000101000)) color_data = 12'b011010011101;
		if(({row_reg, col_reg}==18'b010001000000101001)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b010001000000101010)) color_data = 12'b100110101101;
		if(({row_reg, col_reg}==18'b010001000000101011)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==18'b010001000000101100)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}>=18'b010001000000101101) && ({row_reg, col_reg}<18'b010001000000101111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010001000000101111) && ({row_reg, col_reg}<18'b010001000000111000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001000000111000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010001000000111001) && ({row_reg, col_reg}<18'b010001000000111011)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010001000000111011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010001000000111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010001000000111101)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010001000000111110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010001000000111111)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==18'b010001000001000000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010001000001000001)) color_data = 12'b100010011000;
		if(({row_reg, col_reg}==18'b010001000001000010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010001000001000011)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b010001000001000100)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b010001000001000101)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==18'b010001000001000110)) color_data = 12'b011010001011;
		if(({row_reg, col_reg}==18'b010001000001000111)) color_data = 12'b010101111010;
		if(({row_reg, col_reg}==18'b010001000001001000)) color_data = 12'b010001101010;
		if(({row_reg, col_reg}==18'b010001000001001001)) color_data = 12'b010001101011;
		if(({row_reg, col_reg}==18'b010001000001001010)) color_data = 12'b001101101011;
		if(({row_reg, col_reg}>=18'b010001000001001011) && ({row_reg, col_reg}<18'b010001000001001110)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010001000001001110)) color_data = 12'b001110001011;
		if(({row_reg, col_reg}==18'b010001000001001111)) color_data = 12'b010010001011;
		if(({row_reg, col_reg}==18'b010001000001010000)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}==18'b010001000001010001)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b010001000001010010)) color_data = 12'b101010111100;
		if(({row_reg, col_reg}==18'b010001000001010011)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b010001000001010100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010001000001010101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010001000001010110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010001000001010111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010001000001011000) && ({row_reg, col_reg}<18'b010001000001011100)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010001000001011100) && ({row_reg, col_reg}<18'b010001000001011110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010001000001011110) && ({row_reg, col_reg}<18'b010001000001100000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010001000001100000)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}>=18'b010001000001100001) && ({row_reg, col_reg}<18'b010001000001100011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010001000001100011)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010001000001100100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010001000001100101) && ({row_reg, col_reg}<18'b010001000001100111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010001000001100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010001000001101000) && ({row_reg, col_reg}<18'b010001000001101010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010001000001101010) && ({row_reg, col_reg}<18'b010001000001101100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001000001101100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010001000001101101) && ({row_reg, col_reg}<18'b010001000001101111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010001000001101111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010001000001110000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010001000001110001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010001000001110010) && ({row_reg, col_reg}<18'b010001000001110110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010001000001110110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001000001110111)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b010001000001111000) && ({row_reg, col_reg}<18'b010001000001111100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001000001111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010001000001111101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001000001111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010001000001111111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010001000010000000) && ({row_reg, col_reg}<18'b010001000010000100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b010001000010000100) && ({row_reg, col_reg}<18'b010001000010000111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010001000010000111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010001000010001000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010001000010001001) && ({row_reg, col_reg}<18'b010001000010010011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001000010010011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010001000010010100) && ({row_reg, col_reg}<18'b010001000010010111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b010001000010010111) && ({row_reg, col_reg}<18'b010001000010011100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010001000010011100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010001000010011101) && ({row_reg, col_reg}<18'b010001000010100000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001000010100000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010001000010100001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010001000010100010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010001000010100011)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010001000010100100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010001000010100101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010001000010100110)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==18'b010001000010100111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010001000010101000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b010001000010101001) && ({row_reg, col_reg}<18'b010001000010101011)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010001000010101011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001000010101100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010001000010101101)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b010001000010101110)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==18'b010001000010101111)) color_data = 12'b011010001010;
		if(({row_reg, col_reg}==18'b010001000010110000)) color_data = 12'b010001111010;
		if(({row_reg, col_reg}>=18'b010001000010110001) && ({row_reg, col_reg}<18'b010001000010110011)) color_data = 12'b010101111010;
		if(({row_reg, col_reg}==18'b010001000010110011)) color_data = 12'b011110001010;
		if(({row_reg, col_reg}==18'b010001000010110100)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==18'b010001000010110101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010001000010110110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010001000010110111) && ({row_reg, col_reg}<18'b010001000010111001)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b010001000010111001) && ({row_reg, col_reg}<18'b010001000010111101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010001000010111101)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b010001000010111110) && ({row_reg, col_reg}<18'b010001000011000000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001000011000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010001000011000001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010001000011000010) && ({row_reg, col_reg}<18'b010001000011000100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010001000011000100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010001000011000101) && ({row_reg, col_reg}<18'b010001000011000111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010001000011000111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010001000011001000) && ({row_reg, col_reg}<18'b010001000011001011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010001000011001011)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010001000011001100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==18'b010001000011001101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001000011001110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010001000011001111) && ({row_reg, col_reg}<18'b010001000011010101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b010001000011010101) && ({row_reg, col_reg}<18'b010001000011011000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010001000011011000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001000011011001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010001000011011010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010001000011011011) && ({row_reg, col_reg}<18'b010001000011100011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001000011100011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010001000011100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010001000011100101) && ({row_reg, col_reg}<18'b010001000011101000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010001000011101000) && ({row_reg, col_reg}<18'b010001000011101100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010001000011101100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010001000011101101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001000011101110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010001000011101111) && ({row_reg, col_reg}<18'b010001000011110001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010001000011110001)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}==18'b010001000011110010)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}==18'b010001000011110011)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}==18'b010001000011110100)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}>=18'b010001000011110101) && ({row_reg, col_reg}<18'b010001000011110111)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b010001000011110111)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b010001000011111000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010001000011111001)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}==18'b010001000011111010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010001000011111011)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010001000011111100) && ({row_reg, col_reg}<18'b010001000011111110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010001000011111110) && ({row_reg, col_reg}<18'b010001000100000000)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b010001000100000000) && ({row_reg, col_reg}<18'b010001001000011000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010001001000011000) && ({row_reg, col_reg}<18'b010001001000011011)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010001001000011011) && ({row_reg, col_reg}<18'b010001001000011111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010001001000011111)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010001001000100000) && ({row_reg, col_reg}<18'b010001001000100011)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b010001001000100011)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}==18'b010001001000100100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010001001000100101)) color_data = 12'b010110011101;
		if(({row_reg, col_reg}==18'b010001001000100110)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}==18'b010001001000100111)) color_data = 12'b010010001100;
		if(({row_reg, col_reg}==18'b010001001000101000)) color_data = 12'b010110001100;
		if(({row_reg, col_reg}==18'b010001001000101001)) color_data = 12'b011110011100;
		if(({row_reg, col_reg}==18'b010001001000101010)) color_data = 12'b100110101101;
		if(({row_reg, col_reg}==18'b010001001000101011)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==18'b010001001000101100)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b010001001000101101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010001001000101110) && ({row_reg, col_reg}<18'b010001001000110010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001001000110010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010001001000110011)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b010001001000110100) && ({row_reg, col_reg}<18'b010001001000111001)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b010001001000111001) && ({row_reg, col_reg}<18'b010001001000111011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010001001000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010001001000111100) && ({row_reg, col_reg}<18'b010001001001000000)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010001001001000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010001001001000001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010001001001000010)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==18'b010001001001000011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010001001001000100)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b010001001001000101)) color_data = 12'b101010111100;
		if(({row_reg, col_reg}==18'b010001001001000110)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b010001001001000111)) color_data = 12'b100010011100;
		if(({row_reg, col_reg}==18'b010001001001001000)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==18'b010001001001001001)) color_data = 12'b100010011100;
		if(({row_reg, col_reg}==18'b010001001001001010)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b010001001001001011)) color_data = 12'b100011001111;
		if(({row_reg, col_reg}==18'b010001001001001100)) color_data = 12'b011111001111;
		if(({row_reg, col_reg}>=18'b010001001001001101) && ({row_reg, col_reg}<18'b010001001001001111)) color_data = 12'b011111001110;
		if(({row_reg, col_reg}==18'b010001001001001111)) color_data = 12'b011010111100;
		if(({row_reg, col_reg}==18'b010001001001010000)) color_data = 12'b010110011011;
		if(({row_reg, col_reg}==18'b010001001001010001)) color_data = 12'b011010011011;
		if(({row_reg, col_reg}==18'b010001001001010010)) color_data = 12'b011010001011;
		if(({row_reg, col_reg}==18'b010001001001010011)) color_data = 12'b011010001010;
		if(({row_reg, col_reg}==18'b010001001001010100)) color_data = 12'b100010001010;
		if(({row_reg, col_reg}>=18'b010001001001010101) && ({row_reg, col_reg}<18'b010001001001010111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010001001001010111)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}>=18'b010001001001011000) && ({row_reg, col_reg}<18'b010001001001011011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010001001001011011)) color_data = 12'b100110001001;
		if(({row_reg, col_reg}==18'b010001001001011100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010001001001011101)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010001001001011110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010001001001011111)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==18'b010001001001100000)) color_data = 12'b100001100101;
		if(({row_reg, col_reg}==18'b010001001001100001)) color_data = 12'b100001100110;
		if(({row_reg, col_reg}>=18'b010001001001100010) && ({row_reg, col_reg}<18'b010001001001100100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010001001001100100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010001001001100101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010001001001100110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010001001001100111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001001001101000)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010001001001101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010001001001101010)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010001001001101011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010001001001101100) && ({row_reg, col_reg}<18'b010001001001101110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001001001101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010001001001101111) && ({row_reg, col_reg}<18'b010001001001110001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001001001110001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010001001001110010) && ({row_reg, col_reg}<18'b010001001001110110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010001001001110110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001001001110111)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b010001001001111000) && ({row_reg, col_reg}<18'b010001001001111010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001001001111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010001001001111011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010001001001111100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010001001001111101) && ({row_reg, col_reg}<18'b010001001001111111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010001001001111111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010001001010000000) && ({row_reg, col_reg}<18'b010001001010000100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001001010000100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010001001010000101) && ({row_reg, col_reg}<18'b010001001010001000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010001001010001000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010001001010001001) && ({row_reg, col_reg}<18'b010001001010010011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b010001001010010011) && ({row_reg, col_reg}<18'b010001001010010101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010001001010010101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001001010010110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010001001010010111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b010001001010011000) && ({row_reg, col_reg}<18'b010001001010011100)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010001001010011100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010001001010011101)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010001001010011110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010001001010011111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010001001010100000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001001010100001)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010001001010100010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010001001010100011)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010001001010100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010001001010100101)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010001001010100110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010001001010100111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010001001010101000)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b010001001010101001) && ({row_reg, col_reg}<18'b010001001010101011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010001001010101011) && ({row_reg, col_reg}<18'b010001001010101101)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==18'b010001001010101101)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b010001001010101110)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b010001001010101111)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}==18'b010001001010110000)) color_data = 12'b100010011100;
		if(({row_reg, col_reg}==18'b010001001010110001)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b010001001010110010)) color_data = 12'b100110011100;
		if(({row_reg, col_reg}==18'b010001001010110011)) color_data = 12'b100110011011;
		if(({row_reg, col_reg}==18'b010001001010110100)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}==18'b010001001010110101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010001001010110110)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010001001010110111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010001001010111000) && ({row_reg, col_reg}<18'b010001001010111101)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010001001010111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010001001010111110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001001010111111)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}>=18'b010001001011000000) && ({row_reg, col_reg}<18'b010001001011000010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010001001011000010) && ({row_reg, col_reg}<18'b010001001011000101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010001001011000101) && ({row_reg, col_reg}<18'b010001001011000111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010001001011000111) && ({row_reg, col_reg}<18'b010001001011001011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010001001011001011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010001001011001100) && ({row_reg, col_reg}<18'b010001001011001110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001001011001110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010001001011001111) && ({row_reg, col_reg}<18'b010001001011010101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001001011010101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010001001011010110)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010001001011010111)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==18'b010001001011011000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010001001011011001)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010001001011011010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010001001011011011) && ({row_reg, col_reg}<18'b010001001011100011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001001011100011)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b010001001011100100) && ({row_reg, col_reg}<18'b010001001011101000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010001001011101000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b010001001011101001) && ({row_reg, col_reg}<18'b010001001011101100)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==18'b010001001011101100)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010001001011101101)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010001001011101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010001001011101111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001001011110000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010001001011110001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010001001011110010)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}==18'b010001001011110011)) color_data = 12'b011110001001;
		if(({row_reg, col_reg}==18'b010001001011110100)) color_data = 12'b011110001010;
		if(({row_reg, col_reg}==18'b010001001011110101)) color_data = 12'b011110001011;
		if(({row_reg, col_reg}==18'b010001001011110110)) color_data = 12'b011110011100;
		if(({row_reg, col_reg}==18'b010001001011110111)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b010001001011111000) && ({row_reg, col_reg}<18'b010001001011111010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b010001001011111010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010001001011111011)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010001001011111100) && ({row_reg, col_reg}<18'b010001001011111111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010001001011111111)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b010001001100000000) && ({row_reg, col_reg}<18'b010001010000010111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010001010000010111)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b010001010000011000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010001010000011001) && ({row_reg, col_reg}<18'b010001010000011101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010001010000011101) && ({row_reg, col_reg}<18'b010001010000011111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010001010000011111)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010001010000100000) && ({row_reg, col_reg}<18'b010001010000100010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010001010000100010) && ({row_reg, col_reg}<18'b010001010000100100)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b010001010000100100)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}>=18'b010001010000100101) && ({row_reg, col_reg}<18'b010001010000100111)) color_data = 12'b010001111100;
		if(({row_reg, col_reg}==18'b010001010000100111)) color_data = 12'b010001101011;
		if(({row_reg, col_reg}==18'b010001010000101000)) color_data = 12'b010001111010;
		if(({row_reg, col_reg}==18'b010001010000101001)) color_data = 12'b011010001011;
		if(({row_reg, col_reg}==18'b010001010000101010)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==18'b010001010000101011)) color_data = 12'b101010111100;
		if(({row_reg, col_reg}==18'b010001010000101100)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b010001010000101101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010001010000101110) && ({row_reg, col_reg}<18'b010001010000110011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001010000110011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010001010000110100) && ({row_reg, col_reg}<18'b010001010000111010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010001010000111010) && ({row_reg, col_reg}<18'b010001010000111100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010001010000111100)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}==18'b010001010000111101)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==18'b010001010000111110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010001010000111111)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==18'b010001010001000000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010001010001000001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010001010001000010) && ({row_reg, col_reg}<18'b010001010001000100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001010001000100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010001010001000101)) color_data = 12'b101010111011;
		if(({row_reg, col_reg}>=18'b010001010001000110) && ({row_reg, col_reg}<18'b010001010001001000)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b010001010001001000)) color_data = 12'b101010101100;
		if(({row_reg, col_reg}==18'b010001010001001001)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==18'b010001010001001010)) color_data = 12'b100110111101;
		if(({row_reg, col_reg}==18'b010001010001001011)) color_data = 12'b101011101111;
		if(({row_reg, col_reg}>=18'b010001010001001100) && ({row_reg, col_reg}<18'b010001010001001111)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010001010001001111)) color_data = 12'b100011011110;
		if(({row_reg, col_reg}>=18'b010001010001010000) && ({row_reg, col_reg}<18'b010001010001010010)) color_data = 12'b001101111011;
		if(({row_reg, col_reg}==18'b010001010001010010)) color_data = 12'b001101101011;
		if(({row_reg, col_reg}==18'b010001010001010011)) color_data = 12'b010001101010;
		if(({row_reg, col_reg}==18'b010001010001010100)) color_data = 12'b011110001100;
		if(({row_reg, col_reg}==18'b010001010001010101)) color_data = 12'b101010111100;
		if(({row_reg, col_reg}==18'b010001010001010110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==18'b010001010001010111)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==18'b010001010001011000)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}>=18'b010001010001011001) && ({row_reg, col_reg}<18'b010001010001011011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001010001011011)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==18'b010001010001011100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==18'b010001010001011101)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010001010001011110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010001010001011111) && ({row_reg, col_reg}<18'b010001010001100010)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}>=18'b010001010001100010) && ({row_reg, col_reg}<18'b010001010001100101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010001010001100101)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010001010001100110) && ({row_reg, col_reg}<18'b010001010001101000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010001010001101000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010001010001101001) && ({row_reg, col_reg}<18'b010001010001101100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010001010001101100) && ({row_reg, col_reg}<18'b010001010001110001)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010001010001110001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010001010001110010) && ({row_reg, col_reg}<18'b010001010001110110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010001010001110110) && ({row_reg, col_reg}<18'b010001010001111001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001010001111001)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010001010001111010)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010001010001111011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001010001111100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=18'b010001010001111101) && ({row_reg, col_reg}<18'b010001010010000100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001010010000100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010001010010000101) && ({row_reg, col_reg}<18'b010001010010001000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010001010010001000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010001010010001001) && ({row_reg, col_reg}<18'b010001010010010010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001010010010010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010001010010010011) && ({row_reg, col_reg}<18'b010001010010010101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010001010010010101)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010001010010010110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010001010010010111)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b010001010010011000) && ({row_reg, col_reg}<18'b010001010010011100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001010010011100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010001010010011101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010001010010011110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010001010010011111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010001010010100000)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010001010010100001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010001010010100010)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010001010010100011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010001010010100100) && ({row_reg, col_reg}<18'b010001010010100111)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010001010010100111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010001010010101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010001010010101001) && ({row_reg, col_reg}<18'b010001010010101100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010001010010101100)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==18'b010001010010101101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010001010010101110)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==18'b010001010010101111)) color_data = 12'b101010111011;
		if(({row_reg, col_reg}==18'b010001010010110000)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}>=18'b010001010010110001) && ({row_reg, col_reg}<18'b010001010010110011)) color_data = 12'b101010101100;
		if(({row_reg, col_reg}==18'b010001010010110011)) color_data = 12'b101110101100;
		if(({row_reg, col_reg}>=18'b010001010010110100) && ({row_reg, col_reg}<18'b010001010010110110)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}>=18'b010001010010110110) && ({row_reg, col_reg}<18'b010001010010111010)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010001010010111010)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010001010010111011)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==18'b010001010010111100)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010001010010111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010001010010111110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001010010111111)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}==18'b010001010011000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010001010011000001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001010011000010)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010001010011000011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010001010011000100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010001010011000101) && ({row_reg, col_reg}<18'b010001010011001001)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010001010011001001)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010001010011001010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010001010011001011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010001010011001100) && ({row_reg, col_reg}<18'b010001010011010100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001010011010100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010001010011010101)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b010001010011010110) && ({row_reg, col_reg}<18'b010001010011011001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001010011011001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010001010011011010) && ({row_reg, col_reg}<18'b010001010011100011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001010011100011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010001010011100100) && ({row_reg, col_reg}<18'b010001010011100111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001010011100111)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}>=18'b010001010011101000) && ({row_reg, col_reg}<18'b010001010011101010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b010001010011101010) && ({row_reg, col_reg}<18'b010001010011101100)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==18'b010001010011101100)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010001010011101101)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010001010011101110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001010011101111)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010001010011110000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010001010011110001) && ({row_reg, col_reg}<18'b010001010011110011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010001010011110011)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==18'b010001010011110100)) color_data = 12'b011001111001;
		if(({row_reg, col_reg}==18'b010001010011110101)) color_data = 12'b011001111010;
		if(({row_reg, col_reg}==18'b010001010011110110)) color_data = 12'b011110001011;
		if(({row_reg, col_reg}==18'b010001010011110111)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b010001010011111000) && ({row_reg, col_reg}<18'b010001010011111010)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b010001010011111010) && ({row_reg, col_reg}<18'b010001011000010111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010001011000010111) && ({row_reg, col_reg}<18'b010001011000011011)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010001011000011011) && ({row_reg, col_reg}<18'b010001011000100000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010001011000100000)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==18'b010001011000100001)) color_data = 12'b011010111111;
		if(({row_reg, col_reg}==18'b010001011000100010)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==18'b010001011000100011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010001011000100100)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==18'b010001011000100101)) color_data = 12'b010010001100;
		if(({row_reg, col_reg}>=18'b010001011000100110) && ({row_reg, col_reg}<18'b010001011000101000)) color_data = 12'b010001111011;
		if(({row_reg, col_reg}==18'b010001011000101000)) color_data = 12'b010101111010;
		if(({row_reg, col_reg}==18'b010001011000101001)) color_data = 12'b011110001011;
		if(({row_reg, col_reg}==18'b010001011000101010)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==18'b010001011000101011)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}>=18'b010001011000101100) && ({row_reg, col_reg}<18'b010001011000101110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010001011000101110) && ({row_reg, col_reg}<18'b010001011000110001)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001011000110001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010001011000110010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001011000110011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001011000110100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010001011000110101) && ({row_reg, col_reg}<18'b010001011000110111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010001011000110111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010001011000111000) && ({row_reg, col_reg}<18'b010001011000111010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010001011000111010) && ({row_reg, col_reg}<18'b010001011000111100)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}==18'b010001011000111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010001011000111101)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}>=18'b010001011000111110) && ({row_reg, col_reg}<18'b010001011001000000)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==18'b010001011001000000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010001011001000001) && ({row_reg, col_reg}<18'b010001011001000011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001011001000011)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==18'b010001011001000100)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b010001011001000101) && ({row_reg, col_reg}<18'b010001011001001000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010001011001001000)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==18'b010001011001001001)) color_data = 12'b101010111011;
		if(({row_reg, col_reg}==18'b010001011001001010)) color_data = 12'b100110111011;
		if(({row_reg, col_reg}==18'b010001011001001011)) color_data = 12'b101011101110;
		if(({row_reg, col_reg}>=18'b010001011001001100) && ({row_reg, col_reg}<18'b010001011001001111)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010001011001001111)) color_data = 12'b011111011110;
		if(({row_reg, col_reg}==18'b010001011001010000)) color_data = 12'b001110001011;
		if(({row_reg, col_reg}==18'b010001011001010001)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b010001011001010010)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010001011001010011)) color_data = 12'b001101101100;
		if(({row_reg, col_reg}==18'b010001011001010100)) color_data = 12'b011010011101;
		if(({row_reg, col_reg}==18'b010001011001010101)) color_data = 12'b100110111101;
		if(({row_reg, col_reg}==18'b010001011001010110)) color_data = 12'b101010111011;
		if(({row_reg, col_reg}>=18'b010001011001010111) && ({row_reg, col_reg}<18'b010001011001011010)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b010001011001011010) && ({row_reg, col_reg}<18'b010001011001011100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010001011001011100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==18'b010001011001011101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010001011001011110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010001011001011111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010001011001100000)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==18'b010001011001100001)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}>=18'b010001011001100010) && ({row_reg, col_reg}<18'b010001011001100110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010001011001100110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010001011001100111) && ({row_reg, col_reg}<18'b010001011001110011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010001011001110011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010001011001110100) && ({row_reg, col_reg}<18'b010001011001110110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010001011001110110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001011001110111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010001011001111000) && ({row_reg, col_reg}<18'b010001011001111010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001011001111010)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b010001011001111011) && ({row_reg, col_reg}<18'b010001011001111110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b010001011001111110) && ({row_reg, col_reg}<18'b010001011010000000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010001011010000000) && ({row_reg, col_reg}<18'b010001011010000100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001011010000100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010001011010000101) && ({row_reg, col_reg}<18'b010001011010001000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010001011010001000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010001011010001001) && ({row_reg, col_reg}<18'b010001011010010010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001011010010010)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b010001011010010011) && ({row_reg, col_reg}<18'b010001011010010111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010001011010010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010001011010011000) && ({row_reg, col_reg}<18'b010001011010011100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010001011010011100) && ({row_reg, col_reg}<18'b010001011010011110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010001011010011110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010001011010011111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010001011010100000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001011010100001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010001011010100010) && ({row_reg, col_reg}<18'b010001011010100100)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b010001011010100100) && ({row_reg, col_reg}<18'b010001011010100111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010001011010100111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010001011010101000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010001011010101001) && ({row_reg, col_reg}<18'b010001011010101101)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==18'b010001011010101101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010001011010101110) && ({row_reg, col_reg}<18'b010001011010110000)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}>=18'b010001011010110000) && ({row_reg, col_reg}<18'b010001011010110010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010001011010110010) && ({row_reg, col_reg}<18'b010001011010110100)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==18'b010001011010110100)) color_data = 12'b101010011011;
		if(({row_reg, col_reg}>=18'b010001011010110101) && ({row_reg, col_reg}<18'b010001011010110111)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}>=18'b010001011010110111) && ({row_reg, col_reg}<18'b010001011010111010)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010001011010111010)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==18'b010001011010111011)) color_data = 12'b101010011000;
		if(({row_reg, col_reg}==18'b010001011010111100)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010001011010111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010001011010111110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001011010111111)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}>=18'b010001011011000000) && ({row_reg, col_reg}<18'b010001011011000010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001011011000010)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010001011011000011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010001011011000100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010001011011000101) && ({row_reg, col_reg}<18'b010001011011000111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010001011011000111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010001011011001000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010001011011001001)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010001011011001010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010001011011001011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010001011011001100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010001011011001101) && ({row_reg, col_reg}<18'b010001011011010101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001011011010101)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010001011011010110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001011011010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010001011011011000) && ({row_reg, col_reg}<18'b010001011011100011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001011011100011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010001011011100100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b010001011011100101) && ({row_reg, col_reg}<18'b010001011011100111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010001011011100111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001011011101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010001011011101001) && ({row_reg, col_reg}<18'b010001011011101011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001011011101011)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==18'b010001011011101100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010001011011101101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010001011011101110) && ({row_reg, col_reg}<18'b010001011011110000)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010001011011110000)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010001011011110001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010001011011110010) && ({row_reg, col_reg}<18'b010001011011110100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010001011011110100)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==18'b010001011011110101)) color_data = 12'b011001111001;
		if(({row_reg, col_reg}==18'b010001011011110110)) color_data = 12'b011110001011;
		if(({row_reg, col_reg}==18'b010001011011110111)) color_data = 12'b100010011100;
		if(({row_reg, col_reg}==18'b010001011011111000)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}==18'b010001011011111001)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b010001011011111010) && ({row_reg, col_reg}<18'b010001011011111110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b010001011011111110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010001011011111111)) color_data = 12'b011010101101;

		if(({row_reg, col_reg}>=18'b010001011100000000) && ({row_reg, col_reg}<18'b010001100000011110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010001100000011110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b010001100000011111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010001100000100000)) color_data = 12'b010110101101;
		if(({row_reg, col_reg}==18'b010001100000100001)) color_data = 12'b010110111110;
		if(({row_reg, col_reg}==18'b010001100000100010)) color_data = 12'b010110101101;
		if(({row_reg, col_reg}==18'b010001100000100011)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}==18'b010001100000100100)) color_data = 12'b010110011101;
		if(({row_reg, col_reg}==18'b010001100000100101)) color_data = 12'b010001111011;
		if(({row_reg, col_reg}==18'b010001100000100110)) color_data = 12'b010001101010;
		if(({row_reg, col_reg}==18'b010001100000100111)) color_data = 12'b010101101010;
		if(({row_reg, col_reg}==18'b010001100000101000)) color_data = 12'b010101101001;
		if(({row_reg, col_reg}==18'b010001100000101001)) color_data = 12'b011110001010;
		if(({row_reg, col_reg}==18'b010001100000101010)) color_data = 12'b100110111100;
		if(({row_reg, col_reg}==18'b010001100000101011)) color_data = 12'b101010111011;
		if(({row_reg, col_reg}==18'b010001100000101100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010001100000101101)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}>=18'b010001100000101110) && ({row_reg, col_reg}<18'b010001100000110000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001100000110000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==18'b010001100000110001)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001100000110010)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==18'b010001100000110011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010001100000110100) && ({row_reg, col_reg}<18'b010001100000111001)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010001100000111001)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==18'b010001100000111010)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}==18'b010001100000111011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010001100000111100)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}==18'b010001100000111101)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==18'b010001100000111110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010001100000111111)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}>=18'b010001100001000000) && ({row_reg, col_reg}<18'b010001100001000010)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010001100001000010)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}>=18'b010001100001000011) && ({row_reg, col_reg}<18'b010001100001000101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001100001000101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010001100001000110) && ({row_reg, col_reg}<18'b010001100001001000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b010001100001001000) && ({row_reg, col_reg}<18'b010001100001001010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010001100001001010)) color_data = 12'b100110111011;
		if(({row_reg, col_reg}==18'b010001100001001011)) color_data = 12'b101011101110;
		if(({row_reg, col_reg}==18'b010001100001001100)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010001100001001101) && ({row_reg, col_reg}<18'b010001100001001111)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010001100001001111)) color_data = 12'b011111011110;
		if(({row_reg, col_reg}==18'b010001100001010000)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b010001100001010001)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b010001100001010010)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010001100001010011)) color_data = 12'b010001111101;
		if(({row_reg, col_reg}==18'b010001100001010100)) color_data = 12'b011010011110;
		if(({row_reg, col_reg}==18'b010001100001010101)) color_data = 12'b100010111110;
		if(({row_reg, col_reg}==18'b010001100001010110)) color_data = 12'b100110111101;
		if(({row_reg, col_reg}==18'b010001100001010111)) color_data = 12'b100110111011;
		if(({row_reg, col_reg}>=18'b010001100001011000) && ({row_reg, col_reg}<18'b010001100001011011)) color_data = 12'b101010111011;
		if(({row_reg, col_reg}==18'b010001100001011011)) color_data = 12'b101010111100;
		if(({row_reg, col_reg}==18'b010001100001011100)) color_data = 12'b101010101100;
		if(({row_reg, col_reg}==18'b010001100001011101)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==18'b010001100001011110)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==18'b010001100001011111)) color_data = 12'b010101010101;
		if(({row_reg, col_reg}>=18'b010001100001100000) && ({row_reg, col_reg}<18'b010001100001100010)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==18'b010001100001100010)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010001100001100011) && ({row_reg, col_reg}<18'b010001100001100101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010001100001100101) && ({row_reg, col_reg}<18'b010001100001100111)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==18'b010001100001100111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010001100001101000) && ({row_reg, col_reg}<18'b010001100001110110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010001100001110110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001100001110111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010001100001111000) && ({row_reg, col_reg}<18'b010001100001111010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001100001111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010001100001111011) && ({row_reg, col_reg}<18'b010001100010000100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001100010000100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010001100010000101)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b010001100010000110) && ({row_reg, col_reg}<18'b010001100010001000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010001100010001000)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b010001100010001001) && ({row_reg, col_reg}<18'b010001100010010010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001100010010010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010001100010010011) && ({row_reg, col_reg}<18'b010001100010010111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010001100010010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010001100010011000) && ({row_reg, col_reg}<18'b010001100010011100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001100010011100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010001100010011101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010001100010011110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010001100010011111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010001100010100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010001100010100001)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b010001100010100010) && ({row_reg, col_reg}<18'b010001100010101000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010001100010101000)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010001100010101001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010001100010101010)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==18'b010001100010101011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010001100010101100)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}>=18'b010001100010101101) && ({row_reg, col_reg}<18'b010001100010110000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010001100010110000) && ({row_reg, col_reg}<18'b010001100010110011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001100010110011)) color_data = 12'b101110011010;
		if(({row_reg, col_reg}==18'b010001100010110100)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==18'b010001100010110101)) color_data = 12'b101010011011;
		if(({row_reg, col_reg}>=18'b010001100010110110) && ({row_reg, col_reg}<18'b010001100010111000)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}>=18'b010001100010111000) && ({row_reg, col_reg}<18'b010001100010111011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010001100010111011) && ({row_reg, col_reg}<18'b010001100010111101)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010001100010111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010001100010111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010001100010111111)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}>=18'b010001100011000000) && ({row_reg, col_reg}<18'b010001100011000010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001100011000010)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010001100011000011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010001100011000100) && ({row_reg, col_reg}<18'b010001100011000111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010001100011000111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010001100011001000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010001100011001001)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010001100011001010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010001100011001011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010001100011001100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010001100011001101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001100011001110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010001100011001111) && ({row_reg, col_reg}<18'b010001100011010101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001100011010101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010001100011010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010001100011010111) && ({row_reg, col_reg}<18'b010001100011011101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001100011011101)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b010001100011011110) && ({row_reg, col_reg}<18'b010001100011100011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001100011100011)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}>=18'b010001100011100100) && ({row_reg, col_reg}<18'b010001100011101000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001100011101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010001100011101001)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001100011101010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010001100011101011)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==18'b010001100011101100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010001100011101101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010001100011101110) && ({row_reg, col_reg}<18'b010001100011110000)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010001100011110000) && ({row_reg, col_reg}<18'b010001100011110010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010001100011110010) && ({row_reg, col_reg}<18'b010001100011110100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010001100011110100)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==18'b010001100011110101)) color_data = 12'b011110001001;
		if(({row_reg, col_reg}==18'b010001100011110110)) color_data = 12'b100010011010;
		if(({row_reg, col_reg}==18'b010001100011110111)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}>=18'b010001100011111000) && ({row_reg, col_reg}<18'b010001100011111010)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}>=18'b010001100011111010) && ({row_reg, col_reg}<18'b010001100011111100)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b010001100011111100) && ({row_reg, col_reg}<18'b010001100011111111)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b010001100011111111) && ({row_reg, col_reg}<18'b010001101000010011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010001101000010011) && ({row_reg, col_reg}<18'b010001101000010101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010001101000010101) && ({row_reg, col_reg}<18'b010001101000010111)) color_data = 12'b011110111110;
		if(({row_reg, col_reg}>=18'b010001101000010111) && ({row_reg, col_reg}<18'b010001101000011011)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b010001101000011011)) color_data = 12'b011110111110;
		if(({row_reg, col_reg}==18'b010001101000011100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010001101000011101)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}>=18'b010001101000011110) && ({row_reg, col_reg}<18'b010001101000100000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010001101000100000)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}==18'b010001101000100001)) color_data = 12'b011111001110;
		if(({row_reg, col_reg}==18'b010001101000100010)) color_data = 12'b011011001110;
		if(({row_reg, col_reg}==18'b010001101000100011)) color_data = 12'b011111001111;
		if(({row_reg, col_reg}==18'b010001101000100100)) color_data = 12'b011110111110;
		if(({row_reg, col_reg}==18'b010001101000100101)) color_data = 12'b010110001011;
		if(({row_reg, col_reg}==18'b010001101000100110)) color_data = 12'b011001111011;
		if(({row_reg, col_reg}>=18'b010001101000100111) && ({row_reg, col_reg}<18'b010001101000101001)) color_data = 12'b011001111010;
		if(({row_reg, col_reg}==18'b010001101000101001)) color_data = 12'b100010011010;
		if(({row_reg, col_reg}==18'b010001101000101010)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}>=18'b010001101000101011) && ({row_reg, col_reg}<18'b010001101000101101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010001101000101101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001101000101110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010001101000101111)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}>=18'b010001101000110000) && ({row_reg, col_reg}<18'b010001101000110011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010001101000110011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010001101000110100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010001101000110101) && ({row_reg, col_reg}<18'b010001101000111000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010001101000111000)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010001101000111001) && ({row_reg, col_reg}<18'b010001101000111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010001101000111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010001101000111101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010001101000111110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010001101000111111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010001101001000000)) color_data = 12'b101010011000;
		if(({row_reg, col_reg}==18'b010001101001000001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010001101001000010) && ({row_reg, col_reg}<18'b010001101001001001)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001101001001001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010001101001001010)) color_data = 12'b100110111010;
		if(({row_reg, col_reg}==18'b010001101001001011)) color_data = 12'b101011101110;
		if(({row_reg, col_reg}==18'b010001101001001100)) color_data = 12'b100011111110;
		if(({row_reg, col_reg}==18'b010001101001001101)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010001101001001110)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010001101001001111)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010001101001010000)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b010001101001010001)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010001101001010010)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010001101001010011)) color_data = 12'b010001111101;
		if(({row_reg, col_reg}==18'b010001101001010100)) color_data = 12'b010110001110;
		if(({row_reg, col_reg}==18'b010001101001010101)) color_data = 12'b011110011111;
		if(({row_reg, col_reg}==18'b010001101001010110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b010001101001010111)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b010001101001011000) && ({row_reg, col_reg}<18'b010001101001011010)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b010001101001011010)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}>=18'b010001101001011011) && ({row_reg, col_reg}<18'b010001101001011101)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b010001101001011101)) color_data = 12'b100010011010;
		if(({row_reg, col_reg}==18'b010001101001011110)) color_data = 12'b011110001001;
		if(({row_reg, col_reg}==18'b010001101001011111)) color_data = 12'b011110001000;
		if(({row_reg, col_reg}==18'b010001101001100000)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010001101001100001)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010001101001100010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010001101001100011) && ({row_reg, col_reg}<18'b010001101001100111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010001101001100111)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010001101001101000) && ({row_reg, col_reg}<18'b010001101001110101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010001101001110101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010001101001110110) && ({row_reg, col_reg}<18'b010001101001111010)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010001101001111010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b010001101001111011) && ({row_reg, col_reg}<18'b010001101001111111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b010001101001111111) && ({row_reg, col_reg}<18'b010001101010000101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010001101010000101) && ({row_reg, col_reg}<18'b010001101010000111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010001101010000111) && ({row_reg, col_reg}<18'b010001101010001001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010001101010001001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010001101010001010) && ({row_reg, col_reg}<18'b010001101010001110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b010001101010001110) && ({row_reg, col_reg}<18'b010001101010010000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010001101010010000) && ({row_reg, col_reg}<18'b010001101010010010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001101010010010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010001101010010011) && ({row_reg, col_reg}<18'b010001101010010111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010001101010010111)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b010001101010011000) && ({row_reg, col_reg}<18'b010001101010011100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001101010011100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010001101010011101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010001101010011110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010001101010011111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010001101010100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010001101010100001) && ({row_reg, col_reg}<18'b010001101010100011)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b010001101010100011) && ({row_reg, col_reg}<18'b010001101010100111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010001101010100111) && ({row_reg, col_reg}<18'b010001101010101011)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b010001101010101011) && ({row_reg, col_reg}<18'b010001101010101111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010001101010101111) && ({row_reg, col_reg}<18'b010001101010110001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010001101010110001) && ({row_reg, col_reg}<18'b010001101010110100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001101010110100)) color_data = 12'b100110001001;
		if(({row_reg, col_reg}==18'b010001101010110101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010001101010110110) && ({row_reg, col_reg}<18'b010001101010111000)) color_data = 12'b100110001001;
		if(({row_reg, col_reg}>=18'b010001101010111000) && ({row_reg, col_reg}<18'b010001101010111100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010001101010111100)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010001101010111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010001101010111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010001101010111111) && ({row_reg, col_reg}<18'b010001101011000010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001101011000010)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010001101011000011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010001101011000100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010001101011000101) && ({row_reg, col_reg}<18'b010001101011000111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010001101011000111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001101011001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010001101011001001) && ({row_reg, col_reg}<18'b010001101011001011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001101011001011)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b010001101011001100) && ({row_reg, col_reg}<18'b010001101011010101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001101011010101)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010001101011010110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010001101011010111) && ({row_reg, col_reg}<18'b010001101011011010)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b010001101011011010) && ({row_reg, col_reg}<18'b010001101011011101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001101011011101)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b010001101011011110) && ({row_reg, col_reg}<18'b010001101011100011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001101011100011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010001101011100100)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}>=18'b010001101011100101) && ({row_reg, col_reg}<18'b010001101011101000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001101011101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010001101011101001)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001101011101010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010001101011101011)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==18'b010001101011101100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010001101011101101)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}>=18'b010001101011101110) && ({row_reg, col_reg}<18'b010001101011110000)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010001101011110000)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010001101011110001)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b010001101011110010) && ({row_reg, col_reg}<18'b010001101011110100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001101011110100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010001101011110101)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==18'b010001101011110110)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}==18'b010001101011110111)) color_data = 12'b100010011010;
		if(({row_reg, col_reg}==18'b010001101011111000)) color_data = 12'b100010011011;
		if(({row_reg, col_reg}==18'b010001101011111001)) color_data = 12'b011110011011;
		if(({row_reg, col_reg}==18'b010001101011111010)) color_data = 12'b011110011100;
		if(({row_reg, col_reg}==18'b010001101011111011)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b010001101011111100) && ({row_reg, col_reg}<18'b010001101011111111)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b010001101011111111) && ({row_reg, col_reg}<18'b010001110000001110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010001110000001110) && ({row_reg, col_reg}<18'b010001110000010010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010001110000010010) && ({row_reg, col_reg}<18'b010001110000011100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010001110000011100) && ({row_reg, col_reg}<18'b010001110000011111)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}==18'b010001110000011111)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==18'b010001110000100000)) color_data = 12'b100011011111;
		if(({row_reg, col_reg}>=18'b010001110000100001) && ({row_reg, col_reg}<18'b010001110000100100)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010001110000100100)) color_data = 12'b100111011111;
		if(({row_reg, col_reg}==18'b010001110000100101)) color_data = 12'b100010111101;
		if(({row_reg, col_reg}>=18'b010001110000100110) && ({row_reg, col_reg}<18'b010001110000101000)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==18'b010001110000101000)) color_data = 12'b100110011011;
		if(({row_reg, col_reg}==18'b010001110000101001)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b010001110000101010)) color_data = 12'b101010111011;
		if(({row_reg, col_reg}==18'b010001110000101011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010001110000101100) && ({row_reg, col_reg}<18'b010001110000101110)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==18'b010001110000101110)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010001110000101111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010001110000110000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010001110000110001)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010001110000110010) && ({row_reg, col_reg}<18'b010001110000110101)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010001110000110101) && ({row_reg, col_reg}<18'b010001110000110111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010001110000110111) && ({row_reg, col_reg}<18'b010001110000111011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010001110000111011) && ({row_reg, col_reg}<18'b010001110000111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010001110000111101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001110000111110)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b010001110000111111) && ({row_reg, col_reg}<18'b010001110001000001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001110001000001)) color_data = 12'b101010011000;
		if(({row_reg, col_reg}==18'b010001110001000010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001110001000011)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==18'b010001110001000100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010001110001000101) && ({row_reg, col_reg}<18'b010001110001001001)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001110001001001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010001110001001010)) color_data = 12'b100110111011;
		if(({row_reg, col_reg}==18'b010001110001001011)) color_data = 12'b101011111110;
		if(({row_reg, col_reg}==18'b010001110001001100)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010001110001001101)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010001110001001110)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010001110001001111)) color_data = 12'b100011011111;
		if(({row_reg, col_reg}>=18'b010001110001010000) && ({row_reg, col_reg}<18'b010001110001010010)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010001110001010010)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010001110001010011)) color_data = 12'b001101101100;
		if(({row_reg, col_reg}>=18'b010001110001010100) && ({row_reg, col_reg}<18'b010001110001010111)) color_data = 12'b010001111101;
		if(({row_reg, col_reg}>=18'b010001110001010111) && ({row_reg, col_reg}<18'b010001110001011001)) color_data = 12'b010001111100;
		if(({row_reg, col_reg}>=18'b010001110001011001) && ({row_reg, col_reg}<18'b010001110001011011)) color_data = 12'b010001111011;
		if(({row_reg, col_reg}==18'b010001110001011011)) color_data = 12'b010001111010;
		if(({row_reg, col_reg}==18'b010001110001011100)) color_data = 12'b010001111001;
		if(({row_reg, col_reg}==18'b010001110001011101)) color_data = 12'b011010001010;
		if(({row_reg, col_reg}==18'b010001110001011110)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}==18'b010001110001011111)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}>=18'b010001110001100000) && ({row_reg, col_reg}<18'b010001110001100010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010001110001100010)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010001110001100011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010001110001100100) && ({row_reg, col_reg}<18'b010001110001100110)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010001110001100110) && ({row_reg, col_reg}<18'b010001110001110101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010001110001110101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010001110001110110) && ({row_reg, col_reg}<18'b010001110001111010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010001110001111010) && ({row_reg, col_reg}<18'b010001110001111111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001110001111111)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==18'b010001110010000000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001110010000001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010001110010000010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001110010000011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010001110010000100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010001110010000101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010001110010000110)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b010001110010000111) && ({row_reg, col_reg}<18'b010001110010001001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010001110010001001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010001110010001010) && ({row_reg, col_reg}<18'b010001110010001101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001110010001101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010001110010001110) && ({row_reg, col_reg}<18'b010001110010010000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010001110010010000)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b010001110010010001) && ({row_reg, col_reg}<18'b010001110010010111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010001110010010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010001110010011000) && ({row_reg, col_reg}<18'b010001110010011011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001110010011011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010001110010011100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010001110010011101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010001110010011110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010001110010011111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010001110010100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010001110010100001) && ({row_reg, col_reg}<18'b010001110010100100)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010001110010100100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010001110010100101)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==18'b010001110010100110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010001110010100111)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b010001110010101000) && ({row_reg, col_reg}<18'b010001110010101010)) color_data = 12'b100110101001;
		if(({row_reg, col_reg}>=18'b010001110010101010) && ({row_reg, col_reg}<18'b010001110010101100)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b010001110010101100) && ({row_reg, col_reg}<18'b010001110010101110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010001110010101110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010001110010101111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001110010110000)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}>=18'b010001110010110001) && ({row_reg, col_reg}<18'b010001110010110011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001110010110011)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010001110010110100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010001110010110101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001110010110110)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}==18'b010001110010110111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001110010111000)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010001110010111001)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==18'b010001110010111010)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010001110010111011) && ({row_reg, col_reg}<18'b010001110010111101)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==18'b010001110010111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010001110010111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010001110010111111)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b010001110011000000) && ({row_reg, col_reg}<18'b010001110011000010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010001110011000010) && ({row_reg, col_reg}<18'b010001110011000100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010001110011000100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010001110011000101)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010001110011000110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010001110011000111) && ({row_reg, col_reg}<18'b010001110011001001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010001110011001001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010001110011001010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010001110011001011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010001110011001100) && ({row_reg, col_reg}<18'b010001110011001111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001110011001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010001110011010000) && ({row_reg, col_reg}<18'b010001110011010101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b010001110011010101) && ({row_reg, col_reg}<18'b010001110011010111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010001110011010111) && ({row_reg, col_reg}<18'b010001110011011001)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001110011011001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010001110011011010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010001110011011011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010001110011011100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010001110011011101) && ({row_reg, col_reg}<18'b010001110011011111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010001110011011111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010001110011100000)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010001110011100001) && ({row_reg, col_reg}<18'b010001110011100011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010001110011100011)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b010001110011100100) && ({row_reg, col_reg}<18'b010001110011101010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001110011101010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010001110011101011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b010001110011101100) && ({row_reg, col_reg}<18'b010001110011101111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010001110011101111) && ({row_reg, col_reg}<18'b010001110011110001)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001110011110001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010001110011110010)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b010001110011110011) && ({row_reg, col_reg}<18'b010001110011110101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001110011110101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010001110011110110)) color_data = 12'b011110001000;
		if(({row_reg, col_reg}>=18'b010001110011110111) && ({row_reg, col_reg}<18'b010001110011111001)) color_data = 12'b011110001001;
		if(({row_reg, col_reg}==18'b010001110011111001)) color_data = 12'b011010001001;
		if(({row_reg, col_reg}==18'b010001110011111010)) color_data = 12'b011010001010;
		if(({row_reg, col_reg}==18'b010001110011111011)) color_data = 12'b011110011100;
		if(({row_reg, col_reg}>=18'b010001110011111100) && ({row_reg, col_reg}<18'b010001110011111111)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b010001110011111111) && ({row_reg, col_reg}<18'b010001111000001110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010001111000001110) && ({row_reg, col_reg}<18'b010001111000010001)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010001111000010001) && ({row_reg, col_reg}<18'b010001111000010100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010001111000010100)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}>=18'b010001111000010101) && ({row_reg, col_reg}<18'b010001111000011000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010001111000011000) && ({row_reg, col_reg}<18'b010001111000011011)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b010001111000011011)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}==18'b010001111000011100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010001111000011101)) color_data = 12'b011110111110;
		if(({row_reg, col_reg}==18'b010001111000011110)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}==18'b010001111000011111)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==18'b010001111000100000)) color_data = 12'b100011011111;
		if(({row_reg, col_reg}==18'b010001111000100001)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010001111000100010)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010001111000100011)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b010001111000100100)) color_data = 12'b100111011111;
		if(({row_reg, col_reg}==18'b010001111000100101)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b010001111000100110)) color_data = 12'b100010011100;
		if(({row_reg, col_reg}==18'b010001111000100111)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==18'b010001111000101000)) color_data = 12'b100110011011;
		if(({row_reg, col_reg}==18'b010001111000101001)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}>=18'b010001111000101010) && ({row_reg, col_reg}<18'b010001111000101100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010001111000101100) && ({row_reg, col_reg}<18'b010001111000101110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001111000101110)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010001111000101111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010001111000110000) && ({row_reg, col_reg}<18'b010001111000110010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010001111000110010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010001111000110011) && ({row_reg, col_reg}<18'b010001111000111000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010001111000111000) && ({row_reg, col_reg}<18'b010001111000111010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010001111000111010) && ({row_reg, col_reg}<18'b010001111000111100)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010001111000111100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010001111000111101)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==18'b010001111000111110)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010001111000111111)) color_data = 12'b100010000110;
		if(({row_reg, col_reg}==18'b010001111001000000)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==18'b010001111001000001)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}>=18'b010001111001000010) && ({row_reg, col_reg}<18'b010001111001000101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b010001111001000101) && ({row_reg, col_reg}<18'b010001111001000111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010001111001000111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b010001111001001000) && ({row_reg, col_reg}<18'b010001111001001010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010001111001001010)) color_data = 12'b100010111010;
		if(({row_reg, col_reg}==18'b010001111001001011)) color_data = 12'b100111101101;
		if(({row_reg, col_reg}==18'b010001111001001100)) color_data = 12'b100011111110;
		if(({row_reg, col_reg}>=18'b010001111001001101) && ({row_reg, col_reg}<18'b010001111001001111)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010001111001001111)) color_data = 12'b011111011110;
		if(({row_reg, col_reg}==18'b010001111001010000)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b010001111001010001)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010001111001010010)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}==18'b010001111001010011)) color_data = 12'b010001111101;
		if(({row_reg, col_reg}==18'b010001111001010100)) color_data = 12'b010001111110;
		if(({row_reg, col_reg}==18'b010001111001010101)) color_data = 12'b010001101110;
		if(({row_reg, col_reg}==18'b010001111001010110)) color_data = 12'b001101101110;
		if(({row_reg, col_reg}==18'b010001111001010111)) color_data = 12'b001101101101;
		if(({row_reg, col_reg}==18'b010001111001011000)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b010001111001011001) && ({row_reg, col_reg}<18'b010001111001011011)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010001111001011011)) color_data = 12'b001101111011;
		if(({row_reg, col_reg}==18'b010001111001011100)) color_data = 12'b001101111010;
		if(({row_reg, col_reg}==18'b010001111001011101)) color_data = 12'b010110001010;
		if(({row_reg, col_reg}==18'b010001111001011110)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b010001111001011111)) color_data = 12'b101010111011;
		if(({row_reg, col_reg}==18'b010001111001100000)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==18'b010001111001100001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==18'b010001111001100010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010001111001100011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010001111001100100) && ({row_reg, col_reg}<18'b010001111001100110)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010001111001100110) && ({row_reg, col_reg}<18'b010001111001110101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010001111001110101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010001111001110110) && ({row_reg, col_reg}<18'b010001111001111011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001111001111011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010001111001111100) && ({row_reg, col_reg}<18'b010001111001111111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001111001111111)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b010001111010000000) && ({row_reg, col_reg}<18'b010001111010000100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001111010000100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b010001111010000101) && ({row_reg, col_reg}<18'b010001111010001000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010001111010001000)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b010001111010001001) && ({row_reg, col_reg}<18'b010001111010001101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001111010001101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010001111010001110) && ({row_reg, col_reg}<18'b010001111010010111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010001111010010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010001111010011000) && ({row_reg, col_reg}<18'b010001111010011100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001111010011100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010001111010011101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010001111010011110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010001111010011111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010001111010100000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010001111010100001) && ({row_reg, col_reg}<18'b010001111010100011)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b010001111010100011) && ({row_reg, col_reg}<18'b010001111010100101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010001111010100101) && ({row_reg, col_reg}<18'b010001111010100111)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==18'b010001111010100111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010001111010101000)) color_data = 12'b100110101001;
		if(({row_reg, col_reg}==18'b010001111010101001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010001111010101010)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==18'b010001111010101011)) color_data = 12'b101010101000;
		if(({row_reg, col_reg}==18'b010001111010101100)) color_data = 12'b101010011000;
		if(({row_reg, col_reg}==18'b010001111010101101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010001111010101110)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010001111010101111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010001111010110000)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}>=18'b010001111010110001) && ({row_reg, col_reg}<18'b010001111010110011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001111010110011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010001111010110100) && ({row_reg, col_reg}<18'b010001111010110110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001111010110110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010001111010110111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001111010111000)) color_data = 12'b100110001001;
		if(({row_reg, col_reg}==18'b010001111010111001)) color_data = 12'b101110011010;
		if(({row_reg, col_reg}>=18'b010001111010111010) && ({row_reg, col_reg}<18'b010001111010111101)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==18'b010001111010111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010001111010111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010001111010111111)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b010001111011000000) && ({row_reg, col_reg}<18'b010001111011000010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001111011000010)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010001111011000011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010001111011000100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010001111011000101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010001111011000110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010001111011000111)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b010001111011001000) && ({row_reg, col_reg}<18'b010001111011001010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010001111011001010)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010001111011001011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010001111011001100)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}>=18'b010001111011001101) && ({row_reg, col_reg}<18'b010001111011010011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001111011010011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010001111011010100) && ({row_reg, col_reg}<18'b010001111011010110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001111011010110)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==18'b010001111011010111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==18'b010001111011011000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001111011011001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010001111011011010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010001111011011011) && ({row_reg, col_reg}<18'b010001111011011111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010001111011011111) && ({row_reg, col_reg}<18'b010001111011100011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010001111011100011)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b010001111011100100) && ({row_reg, col_reg}<18'b010001111011101011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b010001111011101011) && ({row_reg, col_reg}<18'b010001111011101101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010001111011101101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010001111011101110)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==18'b010001111011101111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==18'b010001111011110000)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==18'b010001111011110001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010001111011110010) && ({row_reg, col_reg}<18'b010001111011110110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010001111011110110)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==18'b010001111011110111)) color_data = 12'b011110001000;
		if(({row_reg, col_reg}==18'b010001111011111000)) color_data = 12'b011110001001;
		if(({row_reg, col_reg}==18'b010001111011111001)) color_data = 12'b011010001001;
		if(({row_reg, col_reg}==18'b010001111011111010)) color_data = 12'b011010001010;
		if(({row_reg, col_reg}==18'b010001111011111011)) color_data = 12'b011110011100;
		if(({row_reg, col_reg}==18'b010001111011111100)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b010001111011111101) && ({row_reg, col_reg}<18'b010001111011111111)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b010001111011111111) && ({row_reg, col_reg}<18'b010010000000000101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010010000000000101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010010000000000110) && ({row_reg, col_reg}<18'b010010000000001001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010010000000001001)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b010010000000001010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010010000000001011) && ({row_reg, col_reg}<18'b010010000000010000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010010000000010000) && ({row_reg, col_reg}<18'b010010000000010010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010010000000010010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010010000000010011) && ({row_reg, col_reg}<18'b010010000000010101)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}>=18'b010010000000010101) && ({row_reg, col_reg}<18'b010010000000010111)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b010010000000010111)) color_data = 12'b011110111110;
		if(({row_reg, col_reg}==18'b010010000000011000)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b010010000000011001)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}>=18'b010010000000011010) && ({row_reg, col_reg}<18'b010010000000011100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010010000000011100) && ({row_reg, col_reg}<18'b010010000000011110)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==18'b010010000000011110)) color_data = 12'b010110101100;
		if(({row_reg, col_reg}==18'b010010000000011111)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}==18'b010010000000100000)) color_data = 12'b011111101101;
		if(({row_reg, col_reg}>=18'b010010000000100001) && ({row_reg, col_reg}<18'b010010000000100011)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010010000000100011)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}==18'b010010000000100100)) color_data = 12'b101011101110;
		if(({row_reg, col_reg}==18'b010010000000100101)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b010010000000100110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010010000000100111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010010000000101000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b010010000000101001) && ({row_reg, col_reg}<18'b010010000000101011)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010010000000101011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010010000000101100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010010000000101101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010010000000101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010010000000101111)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==18'b010010000000110000)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010010000000110001) && ({row_reg, col_reg}<18'b010010000000110011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010010000000110011) && ({row_reg, col_reg}<18'b010010000000111000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010010000000111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010010000000111001) && ({row_reg, col_reg}<18'b010010000000111011)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010010000000111011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010010000000111100) && ({row_reg, col_reg}<18'b010010000001000000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010000001000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010010000001000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b010010000001000010) && ({row_reg, col_reg}<18'b010010000001000100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b010010000001000100) && ({row_reg, col_reg}<18'b010010000001000110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010010000001000110)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}>=18'b010010000001000111) && ({row_reg, col_reg}<18'b010010000001001001)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==18'b010010000001001001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==18'b010010000001001010)) color_data = 12'b101010111011;
		if(({row_reg, col_reg}==18'b010010000001001011)) color_data = 12'b101011101101;
		if(({row_reg, col_reg}==18'b010010000001001100)) color_data = 12'b101011111110;
		if(({row_reg, col_reg}>=18'b010010000001001101) && ({row_reg, col_reg}<18'b010010000001001111)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010010000001001111)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}==18'b010010000001010000)) color_data = 12'b000110001001;
		if(({row_reg, col_reg}==18'b010010000001010001)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b010010000001010010)) color_data = 12'b000110001100;
		if(({row_reg, col_reg}==18'b010010000001010011)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010010000001010100)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b010010000001010101)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010010000001010110)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}==18'b010010000001010111)) color_data = 12'b001010001110;
		if(({row_reg, col_reg}>=18'b010010000001011000) && ({row_reg, col_reg}<18'b010010000001011010)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010010000001011010)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010010000001011011)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010010000001011100)) color_data = 12'b001101111011;
		if(({row_reg, col_reg}==18'b010010000001011101)) color_data = 12'b010110001011;
		if(({row_reg, col_reg}==18'b010010000001011110)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}==18'b010010000001011111)) color_data = 12'b100110111011;
		if(({row_reg, col_reg}==18'b010010000001100000)) color_data = 12'b100110101001;
		if(({row_reg, col_reg}==18'b010010000001100001)) color_data = 12'b101010111010;
		if(({row_reg, col_reg}==18'b010010000001100010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b010010000001100011) && ({row_reg, col_reg}<18'b010010000001100101)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010010000001100101) && ({row_reg, col_reg}<18'b010010000001100111)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}>=18'b010010000001100111) && ({row_reg, col_reg}<18'b010010000001101100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010010000001101100) && ({row_reg, col_reg}<18'b010010000001101111)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==18'b010010000001101111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010010000001110000) && ({row_reg, col_reg}<18'b010010000001110010)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}>=18'b010010000001110010) && ({row_reg, col_reg}<18'b010010000001110101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010010000001110101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010010000001110110) && ({row_reg, col_reg}<18'b010010000001111111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010010000001111111)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==18'b010010000010000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010010000010000001) && ({row_reg, col_reg}<18'b010010000010000011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010000010000011)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010010000010000100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b010010000010000101) && ({row_reg, col_reg}<18'b010010000010000111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010010000010000111) && ({row_reg, col_reg}<18'b010010000010001001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010010000010001001) && ({row_reg, col_reg}<18'b010010000010001101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010010000010001101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010010000010001110) && ({row_reg, col_reg}<18'b010010000010010011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010010000010010011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010010000010010100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010010000010010101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010010000010010110)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010010000010010111)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b010010000010011000) && ({row_reg, col_reg}<18'b010010000010011100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010000010011100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010010000010011101)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==18'b010010000010011110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010010000010011111)) color_data = 12'b011001010101;
		if(({row_reg, col_reg}==18'b010010000010100000)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010010000010100001) && ({row_reg, col_reg}<18'b010010000010100101)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010010000010100101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010010000010100110)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b010010000010100111) && ({row_reg, col_reg}<18'b010010000010101001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010010000010101001) && ({row_reg, col_reg}<18'b010010000010101011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010010000010101011) && ({row_reg, col_reg}<18'b010010000010101111)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}>=18'b010010000010101111) && ({row_reg, col_reg}<18'b010010000010110001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010010000010110001) && ({row_reg, col_reg}<18'b010010000010110011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010010000010110011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010010000010110100)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010010000010110101)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010010000010110110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010000010110111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010010000010111000)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010010000010111001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010010000010111010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010010000010111011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010010000010111100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010010000010111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010010000010111110) && ({row_reg, col_reg}<18'b010010000011000000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010000011000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010010000011000001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010000011000010)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010010000011000011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010010000011000100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010010000011000101) && ({row_reg, col_reg}<18'b010010000011000111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010010000011000111) && ({row_reg, col_reg}<18'b010010000011001011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010010000011001011)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b010010000011001100) && ({row_reg, col_reg}<18'b010010000011001110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010010000011001110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010010000011001111) && ({row_reg, col_reg}<18'b010010000011011000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b010010000011011000) && ({row_reg, col_reg}<18'b010010000011011010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010010000011011010) && ({row_reg, col_reg}<18'b010010000011011110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010000011011110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010010000011011111) && ({row_reg, col_reg}<18'b010010000011100010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010010000011100010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010010000011100011)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010010000011100100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010010000011100101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010010000011100110) && ({row_reg, col_reg}<18'b010010000011101110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010010000011101110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010010000011101111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010010000011110000)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010010000011110001)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}>=18'b010010000011110010) && ({row_reg, col_reg}<18'b010010000011110111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010010000011110111) && ({row_reg, col_reg}<18'b010010000011111001)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==18'b010010000011111001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010010000011111010)) color_data = 12'b011101111001;
		if(({row_reg, col_reg}==18'b010010000011111011)) color_data = 12'b011110011100;
		if(({row_reg, col_reg}==18'b010010000011111100)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b010010000011111101) && ({row_reg, col_reg}<18'b010010000011111111)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b010010000011111111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010010000100000000)) color_data = 12'b011010101101;

		if(({row_reg, col_reg}>=18'b010010000100000001) && ({row_reg, col_reg}<18'b010010001000000101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010010001000000101) && ({row_reg, col_reg}<18'b010010001000001110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b010010001000001110)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}==18'b010010001000001111)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b010010001000010000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010010001000010001) && ({row_reg, col_reg}<18'b010010001000010011)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b010010001000010011)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}>=18'b010010001000010100) && ({row_reg, col_reg}<18'b010010001000010111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010010001000010111)) color_data = 12'b011110111101;
		if(({row_reg, col_reg}==18'b010010001000011000)) color_data = 12'b011110111110;
		if(({row_reg, col_reg}==18'b010010001000011001)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}==18'b010010001000011010)) color_data = 12'b010110101101;
		if(({row_reg, col_reg}>=18'b010010001000011011) && ({row_reg, col_reg}<18'b010010001000011101)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}==18'b010010001000011101)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}>=18'b010010001000011110) && ({row_reg, col_reg}<18'b010010001000100000)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}==18'b010010001000100000)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}>=18'b010010001000100001) && ({row_reg, col_reg}<18'b010010001000100011)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010010001000100011)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}==18'b010010001000100100)) color_data = 12'b101011011111;
		if(({row_reg, col_reg}==18'b010010001000100101)) color_data = 12'b100110111100;
		if(({row_reg, col_reg}==18'b010010001000100110)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==18'b010010001000100111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010010001000101000) && ({row_reg, col_reg}<18'b010010001000101010)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010010001000101010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010010001000101011) && ({row_reg, col_reg}<18'b010010001000101101)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==18'b010010001000101101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010010001000101110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010010001000101111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010010001000110000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010010001000110001)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}>=18'b010010001000110010) && ({row_reg, col_reg}<18'b010010001000110100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010010001000110100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010010001000110101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010010001000110110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010010001000110111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010010001000111000) && ({row_reg, col_reg}<18'b010010001000111111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010010001000111111) && ({row_reg, col_reg}<18'b010010001001000001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010010001001000001)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}>=18'b010010001001000010) && ({row_reg, col_reg}<18'b010010001001000100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b010010001001000100) && ({row_reg, col_reg}<18'b010010001001001000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010010001001001000)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==18'b010010001001001001)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b010010001001001010)) color_data = 12'b100110111010;
		if(({row_reg, col_reg}==18'b010010001001001011)) color_data = 12'b101111101101;
		if(({row_reg, col_reg}==18'b010010001001001100)) color_data = 12'b101111111110;
		if(({row_reg, col_reg}==18'b010010001001001101)) color_data = 12'b101011111110;
		if(({row_reg, col_reg}==18'b010010001001001110)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b010010001001001111)) color_data = 12'b100011011111;
		if(({row_reg, col_reg}==18'b010010001001010000)) color_data = 12'b001010011010;
		if(({row_reg, col_reg}==18'b010010001001010001)) color_data = 12'b001010001010;
		if(({row_reg, col_reg}==18'b010010001001010010)) color_data = 12'b000101111011;
		if(({row_reg, col_reg}==18'b010010001001010011)) color_data = 12'b001010001101;
		if(({row_reg, col_reg}>=18'b010010001001010100) && ({row_reg, col_reg}<18'b010010001001010111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010010001001010111)) color_data = 12'b001010001101;
		if(({row_reg, col_reg}==18'b010010001001011000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010010001001011001) && ({row_reg, col_reg}<18'b010010001001011011)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010010001001011011)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b010010001001011100)) color_data = 12'b001001111010;
		if(({row_reg, col_reg}==18'b010010001001011101)) color_data = 12'b010010001010;
		if(({row_reg, col_reg}==18'b010010001001011110)) color_data = 12'b011110111100;
		if(({row_reg, col_reg}==18'b010010001001011111)) color_data = 12'b100010111100;
		if(({row_reg, col_reg}==18'b010010001001100000)) color_data = 12'b100110111010;
		if(({row_reg, col_reg}==18'b010010001001100001)) color_data = 12'b101011001011;
		if(({row_reg, col_reg}==18'b010010001001100010)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010010001001100011)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}>=18'b010010001001100100) && ({row_reg, col_reg}<18'b010010001001100110)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==18'b010010001001100110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010010001001100111) && ({row_reg, col_reg}<18'b010010001001110011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010010001001110011)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==18'b010010001001110100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010010001001110101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010010001001110110) && ({row_reg, col_reg}<18'b010010001001111011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010010001001111011)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}>=18'b010010001001111100) && ({row_reg, col_reg}<18'b010010001001111111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010010001001111111)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==18'b010010001010000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010010001010000001) && ({row_reg, col_reg}<18'b010010001010000100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010001010000100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010010001010000101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010010001010000110)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010010001010000111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010010001010001000)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}>=18'b010010001010001001) && ({row_reg, col_reg}<18'b010010001010001011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010010001010001011) && ({row_reg, col_reg}<18'b010010001010001101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010010001010001101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010010001010001110) && ({row_reg, col_reg}<18'b010010001010010000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010010001010010000) && ({row_reg, col_reg}<18'b010010001010010010)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b010010001010010010) && ({row_reg, col_reg}<18'b010010001010010111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010010001010010111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010010001010011000) && ({row_reg, col_reg}<18'b010010001010011100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010001010011100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010010001010011101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010010001010011110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010010001010011111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010010001010100000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010001010100001)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b010010001010100010) && ({row_reg, col_reg}<18'b010010001010100100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010010001010100100)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b010010001010100101) && ({row_reg, col_reg}<18'b010010001010101011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010010001010101011) && ({row_reg, col_reg}<18'b010010001010101110)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==18'b010010001010101110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010010001010101111) && ({row_reg, col_reg}<18'b010010001010110011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010010001010110011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010010001010110100)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b010010001010110101) && ({row_reg, col_reg}<18'b010010001010111000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010001010111000)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010010001010111001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010010001010111010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010010001010111011)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==18'b010010001010111100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010010001010111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010010001010111110) && ({row_reg, col_reg}<18'b010010001011000010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010001011000010)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010010001011000011) && ({row_reg, col_reg}<18'b010010001011000110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010010001011000110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010010001011000111)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b010010001011001000) && ({row_reg, col_reg}<18'b010010001011001010)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010010001011001010)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010010001011001011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010010001011001100) && ({row_reg, col_reg}<18'b010010001011010111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010010001011010111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010010001011011000) && ({row_reg, col_reg}<18'b010010001011011010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010010001011011010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010010001011011011) && ({row_reg, col_reg}<18'b010010001011011110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010001011011110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010010001011011111) && ({row_reg, col_reg}<18'b010010001011100011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010010001011100011)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}>=18'b010010001011100100) && ({row_reg, col_reg}<18'b010010001011101110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b010010001011101110) && ({row_reg, col_reg}<18'b010010001011110000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010010001011110000)) color_data = 12'b101010111010;
		if(({row_reg, col_reg}==18'b010010001011110001)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010010001011110010)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b010010001011110011) && ({row_reg, col_reg}<18'b010010001011110101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010001011110101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010010001011110110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010001011110111)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==18'b010010001011111000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010001011111001)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==18'b010010001011111010)) color_data = 12'b011001111000;
		if(({row_reg, col_reg}==18'b010010001011111011)) color_data = 12'b011110011100;
		if(({row_reg, col_reg}==18'b010010001011111100)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b010010001011111101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010010001011111110) && ({row_reg, col_reg}<18'b010010001100000000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010010001100000000)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b010010001100000001) && ({row_reg, col_reg}<18'b010010010000000100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010010010000000100) && ({row_reg, col_reg}<18'b010010010000001011)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b010010010000001011)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}>=18'b010010010000001100) && ({row_reg, col_reg}<18'b010010010000001110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b010010010000001110)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}>=18'b010010010000001111) && ({row_reg, col_reg}<18'b010010010000010001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010010010000010001)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}==18'b010010010000010010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010010010000010011)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010010010000010100) && ({row_reg, col_reg}<18'b010010010000010110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010010010000010110)) color_data = 12'b011111001111;
		if(({row_reg, col_reg}>=18'b010010010000010111) && ({row_reg, col_reg}<18'b010010010000011001)) color_data = 12'b100011011111;
		if(({row_reg, col_reg}==18'b010010010000011001)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}>=18'b010010010000011010) && ({row_reg, col_reg}<18'b010010010000011111)) color_data = 12'b100011011111;
		if(({row_reg, col_reg}==18'b010010010000011111)) color_data = 12'b011111011110;
		if(({row_reg, col_reg}==18'b010010010000100000)) color_data = 12'b010111001110;
		if(({row_reg, col_reg}==18'b010010010000100001)) color_data = 12'b010110111101;
		if(({row_reg, col_reg}==18'b010010010000100010)) color_data = 12'b010010101100;
		if(({row_reg, col_reg}==18'b010010010000100011)) color_data = 12'b010110101101;
		if(({row_reg, col_reg}==18'b010010010000100100)) color_data = 12'b011010101100;
		if(({row_reg, col_reg}==18'b010010010000100101)) color_data = 12'b011010001001;
		if(({row_reg, col_reg}==18'b010010010000100110)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==18'b010010010000100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010010010000101000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010010010000101001) && ({row_reg, col_reg}<18'b010010010000101011)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010010010000101011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010010000101100)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010010010000101101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010010010000101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010010010000101111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010010010000110000)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010010010000110001)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010010010000110010) && ({row_reg, col_reg}<18'b010010010000110111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010010010000110111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010010010000111000) && ({row_reg, col_reg}<18'b010010010000111100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010010000111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010010010000111101) && ({row_reg, col_reg}<18'b010010010000111111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010010010000111111) && ({row_reg, col_reg}<18'b010010010001000001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010010010001000001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010010010001000010) && ({row_reg, col_reg}<18'b010010010001000100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b010010010001000100) && ({row_reg, col_reg}<18'b010010010001000110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010010010001000110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b010010010001000111) && ({row_reg, col_reg}<18'b010010010001001001)) color_data = 12'b100110001001;
		if(({row_reg, col_reg}==18'b010010010001001001)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010010010001001010)) color_data = 12'b100010011000;
		if(({row_reg, col_reg}==18'b010010010001001011)) color_data = 12'b100010101001;
		if(({row_reg, col_reg}==18'b010010010001001100)) color_data = 12'b100010101010;
		if(({row_reg, col_reg}==18'b010010010001001101)) color_data = 12'b011110101010;
		if(({row_reg, col_reg}==18'b010010010001001110)) color_data = 12'b011110111100;
		if(({row_reg, col_reg}==18'b010010010001001111)) color_data = 12'b100011001101;
		if(({row_reg, col_reg}==18'b010010010001010000)) color_data = 12'b010110111100;
		if(({row_reg, col_reg}==18'b010010010001010001)) color_data = 12'b011011011110;
		if(({row_reg, col_reg}==18'b010010010001010010)) color_data = 12'b011011011111;
		if(({row_reg, col_reg}==18'b010010010001010011)) color_data = 12'b011011001111;
		if(({row_reg, col_reg}==18'b010010010001010100)) color_data = 12'b010110101110;
		if(({row_reg, col_reg}==18'b010010010001010101)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b010010010001010110)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010010010001010111)) color_data = 12'b001010001101;
		if(({row_reg, col_reg}==18'b010010010001011000)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b010010010001011001)) color_data = 12'b010110101110;
		if(({row_reg, col_reg}>=18'b010010010001011010) && ({row_reg, col_reg}<18'b010010010001011100)) color_data = 12'b011111001111;
		if(({row_reg, col_reg}==18'b010010010001011100)) color_data = 12'b011011001110;
		if(({row_reg, col_reg}==18'b010010010001011101)) color_data = 12'b011111001101;
		if(({row_reg, col_reg}>=18'b010010010001011110) && ({row_reg, col_reg}<18'b010010010001100000)) color_data = 12'b100011011110;
		if(({row_reg, col_reg}==18'b010010010001100000)) color_data = 12'b100111001100;
		if(({row_reg, col_reg}==18'b010010010001100001)) color_data = 12'b101011011100;
		if(({row_reg, col_reg}==18'b010010010001100010)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==18'b010010010001100011)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}==18'b010010010001100100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010010010001100101) && ({row_reg, col_reg}<18'b010010010001110010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010010010001110010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010010010001110011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010010010001110100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010010010001110101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010010010001110110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010010010001110111) && ({row_reg, col_reg}<18'b010010010001111011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010010010001111011)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}>=18'b010010010001111100) && ({row_reg, col_reg}<18'b010010010001111111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010010010001111111)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}>=18'b010010010010000000) && ({row_reg, col_reg}<18'b010010010010000100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010010010000100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b010010010010000101) && ({row_reg, col_reg}<18'b010010010010001000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010010010010001000) && ({row_reg, col_reg}<18'b010010010010001011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010010010010001011) && ({row_reg, col_reg}<18'b010010010010001101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010010010010001101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010010010010001110) && ({row_reg, col_reg}<18'b010010010010010010)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010010010010010010) && ({row_reg, col_reg}<18'b010010010010010111)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010010010010010111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010010010011000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010010010010011001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010010010010011010) && ({row_reg, col_reg}<18'b010010010010011101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010010010011101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010010010010011110) && ({row_reg, col_reg}<18'b010010010010100000)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010010010010100000)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==18'b010010010010100001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010010010010100010) && ({row_reg, col_reg}<18'b010010010010100101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010010010010100101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b010010010010100110) && ({row_reg, col_reg}<18'b010010010010110000)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010010010010110000)) color_data = 12'b100110001001;
		if(({row_reg, col_reg}>=18'b010010010010110001) && ({row_reg, col_reg}<18'b010010010010110100)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==18'b010010010010110100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010010010010110101) && ({row_reg, col_reg}<18'b010010010010110111)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==18'b010010010010110111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010010010010111000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b010010010010111001) && ({row_reg, col_reg}<18'b010010010010111101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010010010010111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010010010010111110) && ({row_reg, col_reg}<18'b010010010011000010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010010011000010)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010010010011000011) && ({row_reg, col_reg}<18'b010010010011000110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010010010011000110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010010010011000111) && ({row_reg, col_reg}<18'b010010010011001011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010010010011001011) && ({row_reg, col_reg}<18'b010010010011011010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b010010010011011010) && ({row_reg, col_reg}<18'b010010010011011100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b010010010011011100) && ({row_reg, col_reg}<18'b010010010011011110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010010010011011110) && ({row_reg, col_reg}<18'b010010010011100000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010010010011100000)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==18'b010010010011100001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010010010011100010)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010010010011100011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010010010011100100) && ({row_reg, col_reg}<18'b010010010011101010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b010010010011101010) && ({row_reg, col_reg}<18'b010010010011101100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010010010011101100) && ({row_reg, col_reg}<18'b010010010011101110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010010010011101110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010010010011101111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010010010011110000)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==18'b010010010011110001)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010010010011110010)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==18'b010010010011110011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b010010010011110100) && ({row_reg, col_reg}<18'b010010010011110110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010010010011110110)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010010010011110111)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010010010011111000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010010011111001)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==18'b010010010011111010)) color_data = 12'b011110001001;
		if(({row_reg, col_reg}==18'b010010010011111011)) color_data = 12'b011110011100;
		if(({row_reg, col_reg}==18'b010010010011111100)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b010010010011111101) && ({row_reg, col_reg}<18'b010010010011111111)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010010010011111111) && ({row_reg, col_reg}<18'b010010010100000100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010010010100000100)) color_data = 12'b011010101111;

		if(({row_reg, col_reg}>=18'b010010010100000101) && ({row_reg, col_reg}<18'b010010011000000000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010010011000000000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b010010011000000001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010010011000000010) && ({row_reg, col_reg}<18'b010010011000000101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b010010011000000101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010010011000000110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010010011000000111) && ({row_reg, col_reg}<18'b010010011000001001)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}==18'b010010011000001001)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b010010011000001010)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}==18'b010010011000001011)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010010011000001100) && ({row_reg, col_reg}<18'b010010011000001110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010010011000001110) && ({row_reg, col_reg}<18'b010010011000010000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b010010011000010000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010010011000010001)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}==18'b010010011000010010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010010011000010011) && ({row_reg, col_reg}<18'b010010011000010101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010010011000010101)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==18'b010010011000010110)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}>=18'b010010011000010111) && ({row_reg, col_reg}<18'b010010011000011010)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010010011000011010)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010010011000011011) && ({row_reg, col_reg}<18'b010010011000011110)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010010011000011110)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}==18'b010010011000011111)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010010011000100000)) color_data = 12'b001110011100;
		if(({row_reg, col_reg}==18'b010010011000100001)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}>=18'b010010011000100010) && ({row_reg, col_reg}<18'b010010011000100100)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b010010011000100100)) color_data = 12'b001101101010;
		if(({row_reg, col_reg}==18'b010010011000100101)) color_data = 12'b010101111001;
		if(({row_reg, col_reg}==18'b010010011000100110)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}==18'b010010011000100111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010010011000101000) && ({row_reg, col_reg}<18'b010010011000101010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010010011000101010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010010011000101011) && ({row_reg, col_reg}<18'b010010011000101110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010010011000101110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010010011000101111)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}==18'b010010011000110000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010010011000110001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010010011000110010)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010010011000110011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010011000110100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010010011000110101)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b010010011000110110) && ({row_reg, col_reg}<18'b010010011000111100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010011000111100)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b010010011000111101) && ({row_reg, col_reg}<18'b010010011001000000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010010011001000000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=18'b010010011001000001) && ({row_reg, col_reg}<18'b010010011001000100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b010010011001000100) && ({row_reg, col_reg}<18'b010010011001000110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010010011001000110)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010010011001000111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010011001001000)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}>=18'b010010011001001001) && ({row_reg, col_reg}<18'b010010011001001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010010011001001011) && ({row_reg, col_reg}<18'b010010011001001101)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==18'b010010011001001101)) color_data = 12'b011010001000;
		if(({row_reg, col_reg}==18'b010010011001001110)) color_data = 12'b011010001001;
		if(({row_reg, col_reg}==18'b010010011001001111)) color_data = 12'b011010011010;
		if(({row_reg, col_reg}==18'b010010011001010000)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}>=18'b010010011001010001) && ({row_reg, col_reg}<18'b010010011001010100)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010010011001010100)) color_data = 12'b011011001110;
		if(({row_reg, col_reg}==18'b010010011001010101)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}>=18'b010010011001010110) && ({row_reg, col_reg}<18'b010010011001011001)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b010010011001011001)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}>=18'b010010011001011010) && ({row_reg, col_reg}<18'b010010011001011100)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010010011001011100)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}>=18'b010010011001011101) && ({row_reg, col_reg}<18'b010010011001100000)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010010011001100000)) color_data = 12'b101011111110;
		if(({row_reg, col_reg}==18'b010010011001100001)) color_data = 12'b101111101110;
		if(({row_reg, col_reg}==18'b010010011001100010)) color_data = 12'b101011001100;
		if(({row_reg, col_reg}==18'b010010011001100011)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==18'b010010011001100100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010010011001100101) && ({row_reg, col_reg}<18'b010010011001101010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010010011001101010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010010011001101011) && ({row_reg, col_reg}<18'b010010011001101101)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}>=18'b010010011001101101) && ({row_reg, col_reg}<18'b010010011001110000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010010011001110000) && ({row_reg, col_reg}<18'b010010011001110011)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==18'b010010011001110011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010010011001110100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010010011001110101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010010011001110110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010010011001110111) && ({row_reg, col_reg}<18'b010010011001111111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010010011001111111)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010010011010000000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010011010000001)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}>=18'b010010011010000010) && ({row_reg, col_reg}<18'b010010011010000100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010011010000100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010010011010000101) && ({row_reg, col_reg}<18'b010010011010000111)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010010011010000111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010010011010001000)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010010011010001001)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==18'b010010011010001010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b010010011010001011) && ({row_reg, col_reg}<18'b010010011010001110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010010011010001110)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b010010011010001111) && ({row_reg, col_reg}<18'b010010011010010010)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010010011010010010)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b010010011010010011) && ({row_reg, col_reg}<18'b010010011010010111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010011010010111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010010011010011000) && ({row_reg, col_reg}<18'b010010011010011011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010010011010011011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010010011010011100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010010011010011101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010010011010011110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010010011010011111) && ({row_reg, col_reg}<18'b010010011010100001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010010011010100001)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b010010011010100010) && ({row_reg, col_reg}<18'b010010011010100101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010010011010100101)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b010010011010100110) && ({row_reg, col_reg}<18'b010010011010110011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010011010110011)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b010010011010110100) && ({row_reg, col_reg}<18'b010010011010110110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010010011010110110)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010010011010110111)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==18'b010010011010111000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010010011010111001) && ({row_reg, col_reg}<18'b010010011010111101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010010011010111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010010011010111110) && ({row_reg, col_reg}<18'b010010011011000010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010011011000010)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010010011011000011) && ({row_reg, col_reg}<18'b010010011011000110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010010011011000110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010010011011000111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010010011011001000) && ({row_reg, col_reg}<18'b010010011011011010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010010011011011010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010010011011011011) && ({row_reg, col_reg}<18'b010010011011100110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010010011011100110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010010011011100111) && ({row_reg, col_reg}<18'b010010011011110100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010010011011110100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==18'b010010011011110101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010010011011110110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010010011011110111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010010011011111000) && ({row_reg, col_reg}<18'b010010011011111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010010011011111010)) color_data = 12'b011110001001;
		if(({row_reg, col_reg}==18'b010010011011111011)) color_data = 12'b011110011011;
		if(({row_reg, col_reg}==18'b010010011011111100)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b010010011011111101) && ({row_reg, col_reg}<18'b010010011011111111)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010010011011111111) && ({row_reg, col_reg}<18'b010010011100000011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010010011100000011) && ({row_reg, col_reg}<18'b010010011100000110)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b010010011100000110) && ({row_reg, col_reg}<18'b010010011100001001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010010011100001001)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b010010011100001010) && ({row_reg, col_reg}<18'b010010100000000010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010010100000000010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b010010100000000011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010010100000000100)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010010100000000101) && ({row_reg, col_reg}<18'b010010100000001110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010010100000001110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b010010100000001111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010010100000010000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b010010100000010001)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}==18'b010010100000010010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010010100000010011) && ({row_reg, col_reg}<18'b010010100000010101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010010100000010101)) color_data = 12'b010110101101;
		if(({row_reg, col_reg}==18'b010010100000010110)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}==18'b010010100000010111)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010010100000011000) && ({row_reg, col_reg}<18'b010010100000011101)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010010100000011101)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010010100000011110)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010010100000011111)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b010010100000100000)) color_data = 12'b001110011101;
		if(({row_reg, col_reg}==18'b010010100000100001)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b010010100000100010) && ({row_reg, col_reg}<18'b010010100000100100)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b010010100000100100)) color_data = 12'b010001111011;
		if(({row_reg, col_reg}==18'b010010100000100101)) color_data = 12'b010101111001;
		if(({row_reg, col_reg}==18'b010010100000100110)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}==18'b010010100000100111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010010100000101000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010010100000101001)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010010100000101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010010100000101011)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010010100000101100) && ({row_reg, col_reg}<18'b010010100000101111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010010100000101111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010010100000110000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010010100000110001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010010100000110010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010010100000110011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010010100000110100) && ({row_reg, col_reg}<18'b010010100000111001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010100000111001)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b010010100000111010) && ({row_reg, col_reg}<18'b010010100000111100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010100000111100)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b010010100000111101) && ({row_reg, col_reg}<18'b010010100000111111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010010100000111111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010010100001000000) && ({row_reg, col_reg}<18'b010010100001000010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b010010100001000010) && ({row_reg, col_reg}<18'b010010100001000100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010010100001000100)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010010100001000101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010010100001000110)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010010100001000111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010100001001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010010100001001001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010010100001001010) && ({row_reg, col_reg}<18'b010010100001001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010010100001001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010010100001001101)) color_data = 12'b011110001000;
		if(({row_reg, col_reg}==18'b010010100001001110)) color_data = 12'b011001111000;
		if(({row_reg, col_reg}==18'b010010100001001111)) color_data = 12'b011110011010;
		if(({row_reg, col_reg}==18'b010010100001010000)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}==18'b010010100001010001)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b010010100001010010)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010010100001010011)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010010100001010100)) color_data = 12'b010110111101;
		if(({row_reg, col_reg}==18'b010010100001010101)) color_data = 12'b000101111010;
		if(({row_reg, col_reg}==18'b010010100001010110)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b010010100001010111)) color_data = 12'b001010001101;
		if(({row_reg, col_reg}==18'b010010100001011000)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b010010100001011001)) color_data = 12'b011111001111;
		if(({row_reg, col_reg}>=18'b010010100001011010) && ({row_reg, col_reg}<18'b010010100001011101)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010010100001011101) && ({row_reg, col_reg}<18'b010010100001100000)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010010100001100000)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}==18'b010010100001100001)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b010010100001100010)) color_data = 12'b100111011101;
		if(({row_reg, col_reg}==18'b010010100001100011)) color_data = 12'b010101110111;
		if(({row_reg, col_reg}==18'b010010100001100100)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==18'b010010100001100101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010010100001100110) && ({row_reg, col_reg}<18'b010010100001101010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010010100001101010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010010100001101011) && ({row_reg, col_reg}<18'b010010100001101101)) color_data = 12'b011001110101;
		if(({row_reg, col_reg}==18'b010010100001101101)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}>=18'b010010100001101110) && ({row_reg, col_reg}<18'b010010100001110000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010010100001110000) && ({row_reg, col_reg}<18'b010010100001110010)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==18'b010010100001110010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010010100001110011)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010010100001110100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010010100001110101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010010100001110110)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010010100001110111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010010100001111000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010010100001111001)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010010100001111010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010010100001111011) && ({row_reg, col_reg}<18'b010010100001111110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010010100001111110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010010100001111111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010010100010000000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010100010000001)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==18'b010010100010000010)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010010100010000011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010100010000100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010010100010000101) && ({row_reg, col_reg}<18'b010010100010000111)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010010100010000111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010010100010001000)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010010100010001001)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}>=18'b010010100010001010) && ({row_reg, col_reg}<18'b010010100010001100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b010010100010001100) && ({row_reg, col_reg}<18'b010010100010001110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010010100010001110)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010010100010001111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010010100010010000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010010100010010001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010010100010010010)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b010010100010010011) && ({row_reg, col_reg}<18'b010010100010010111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010100010010111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010010100010011000) && ({row_reg, col_reg}<18'b010010100010011011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010010100010011011)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010010100010011100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010010100010011101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010010100010011110) && ({row_reg, col_reg}<18'b010010100010100100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010010100010100100)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010010100010100101)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}>=18'b010010100010100110) && ({row_reg, col_reg}<18'b010010100010110011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010100010110011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010010100010110100) && ({row_reg, col_reg}<18'b010010100010110110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010010100010110110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010010100010110111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b010010100010111000) && ({row_reg, col_reg}<18'b010010100010111010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010010100010111010) && ({row_reg, col_reg}<18'b010010100010111100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010010100010111100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010010100010111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010010100010111110) && ({row_reg, col_reg}<18'b010010100011000010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010100011000010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010010100011000011) && ({row_reg, col_reg}<18'b010010100011000110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010010100011000110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010010100011000111) && ({row_reg, col_reg}<18'b010010100011100100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010010100011100100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==18'b010010100011100101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010010100011100110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010010100011100111) && ({row_reg, col_reg}<18'b010010100011101001)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010010100011101001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010010100011101010) && ({row_reg, col_reg}<18'b010010100011110000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b010010100011110000) && ({row_reg, col_reg}<18'b010010100011110010)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==18'b010010100011110010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010010100011110011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010010100011110100) && ({row_reg, col_reg}<18'b010010100011110110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010010100011110110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010010100011110111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010010100011111000) && ({row_reg, col_reg}<18'b010010100011111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010010100011111010)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==18'b010010100011111011)) color_data = 12'b011110011011;
		if(({row_reg, col_reg}==18'b010010100011111100)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}==18'b010010100011111101)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b010010100011111110) && ({row_reg, col_reg}<18'b010010100100000010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b010010100100000010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010010100100000011) && ({row_reg, col_reg}<18'b010010100100000101)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b010010100100000101) && ({row_reg, col_reg}<18'b010010100100001001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010010100100001001)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b010010100100001010) && ({row_reg, col_reg}<18'b010010101000000100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010010101000000100)) color_data = 12'b011110111110;
		if(({row_reg, col_reg}>=18'b010010101000000101) && ({row_reg, col_reg}<18'b010010101000000111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010010101000000111) && ({row_reg, col_reg}<18'b010010101000001001)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}>=18'b010010101000001001) && ({row_reg, col_reg}<18'b010010101000001101)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}>=18'b010010101000001101) && ({row_reg, col_reg}<18'b010010101000001111)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}==18'b010010101000001111)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}==18'b010010101000010000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010010101000010001)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b010010101000010010)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}==18'b010010101000010011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010010101000010100)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}==18'b010010101000010101)) color_data = 12'b010110101101;
		if(({row_reg, col_reg}==18'b010010101000010110)) color_data = 12'b011111011110;
		if(({row_reg, col_reg}==18'b010010101000010111)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010010101000011000) && ({row_reg, col_reg}<18'b010010101000011011)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010010101000011011)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010010101000011100) && ({row_reg, col_reg}<18'b010010101000011110)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010010101000011110)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010010101000011111)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010010101000100000)) color_data = 12'b001110011101;
		if(({row_reg, col_reg}==18'b010010101000100001)) color_data = 12'b000101111011;
		if(({row_reg, col_reg}==18'b010010101000100010)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b010010101000100011)) color_data = 12'b001101111011;
		if(({row_reg, col_reg}==18'b010010101000100100)) color_data = 12'b010001111010;
		if(({row_reg, col_reg}==18'b010010101000100101)) color_data = 12'b010101101000;
		if(({row_reg, col_reg}==18'b010010101000100110)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010010101000100111) && ({row_reg, col_reg}<18'b010010101000101011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010010101000101011)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010010101000101100) && ({row_reg, col_reg}<18'b010010101000101111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010010101000101111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010010101000110000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010010101000110001) && ({row_reg, col_reg}<18'b010010101000110011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010010101000110011) && ({row_reg, col_reg}<18'b010010101000110101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010010101000110101) && ({row_reg, col_reg}<18'b010010101000111010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010010101000111010) && ({row_reg, col_reg}<18'b010010101000111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010010101000111100)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b010010101000111101) && ({row_reg, col_reg}<18'b010010101000111111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010010101000111111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010010101001000000) && ({row_reg, col_reg}<18'b010010101001000101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010010101001000101)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==18'b010010101001000110)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b010010101001000111) && ({row_reg, col_reg}<18'b010010101001001001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010101001001001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010010101001001010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010101001001011)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010010101001001100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010101001001101)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}==18'b010010101001001110)) color_data = 12'b011110001000;
		if(({row_reg, col_reg}==18'b010010101001001111)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}==18'b010010101001010000)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}==18'b010010101001010001)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}>=18'b010010101001010010) && ({row_reg, col_reg}<18'b010010101001010100)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010010101001010100)) color_data = 12'b010110111110;
		if(({row_reg, col_reg}==18'b010010101001010101)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b010010101001010110)) color_data = 12'b001010001101;
		if(({row_reg, col_reg}==18'b010010101001010111)) color_data = 12'b001010001110;
		if(({row_reg, col_reg}==18'b010010101001011000)) color_data = 12'b001010001101;
		if(({row_reg, col_reg}==18'b010010101001011001)) color_data = 12'b011111001111;
		if(({row_reg, col_reg}==18'b010010101001011010)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}>=18'b010010101001011011) && ({row_reg, col_reg}<18'b010010101001011101)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010010101001011101) && ({row_reg, col_reg}<18'b010010101001100000)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010010101001100000) && ({row_reg, col_reg}<18'b010010101001100010)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010010101001100010)) color_data = 12'b100111011110;
		if(({row_reg, col_reg}==18'b010010101001100011)) color_data = 12'b010001111000;
		if(({row_reg, col_reg}==18'b010010101001100100)) color_data = 12'b010101110111;
		if(({row_reg, col_reg}==18'b010010101001100101)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==18'b010010101001100110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010010101001100111) && ({row_reg, col_reg}<18'b010010101001101011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010010101001101011)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==18'b010010101001101100)) color_data = 12'b011001110101;
		if(({row_reg, col_reg}==18'b010010101001101101)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}>=18'b010010101001101110) && ({row_reg, col_reg}<18'b010010101001110000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010010101001110000)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010010101001110001) && ({row_reg, col_reg}<18'b010010101001110011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010010101001110011)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010010101001110100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010010101001110101)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010010101001110110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010010101001110111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b010010101001111000) && ({row_reg, col_reg}<18'b010010101001111011)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==18'b010010101001111011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=18'b010010101001111100) && ({row_reg, col_reg}<18'b010010101001111111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010010101001111111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010010101010000000)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010010101010000001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010101010000010)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010010101010000011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010101010000100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010010101010000101) && ({row_reg, col_reg}<18'b010010101010000111)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010010101010000111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010010101010001000)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b010010101010001001) && ({row_reg, col_reg}<18'b010010101010001101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b010010101010001101) && ({row_reg, col_reg}<18'b010010101010001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010010101010001111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010010101010010000)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010010101010010001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010010101010010010)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b010010101010010011) && ({row_reg, col_reg}<18'b010010101010010111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010101010010111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010010101010011000) && ({row_reg, col_reg}<18'b010010101010011011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010010101010011011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010101010011100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010010101010011101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010010101010011110) && ({row_reg, col_reg}<18'b010010101010100000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010010101010100000)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010010101010100001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010010101010100010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010010101010100011) && ({row_reg, col_reg}<18'b010010101010100101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010010101010100101)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b010010101010100110) && ({row_reg, col_reg}<18'b010010101010110011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010101010110011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010010101010110100) && ({row_reg, col_reg}<18'b010010101010111000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010010101010111000)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010010101010111001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010010101010111010) && ({row_reg, col_reg}<18'b010010101010111100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010010101010111100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010010101010111101)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b010010101010111110) && ({row_reg, col_reg}<18'b010010101011000010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010101011000010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010010101011000011) && ({row_reg, col_reg}<18'b010010101011000110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010010101011000110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010010101011000111) && ({row_reg, col_reg}<18'b010010101011101110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b010010101011101110) && ({row_reg, col_reg}<18'b010010101011110001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010010101011110001) && ({row_reg, col_reg}<18'b010010101011110100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010010101011110100)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==18'b010010101011110101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010010101011110110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010010101011110111)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b010010101011111000) && ({row_reg, col_reg}<18'b010010101011111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010010101011111010)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==18'b010010101011111011)) color_data = 12'b100010011011;
		if(({row_reg, col_reg}==18'b010010101011111100)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}>=18'b010010101011111101) && ({row_reg, col_reg}<18'b010010101100000000)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b010010101100000000) && ({row_reg, col_reg}<18'b010010101100000010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010010101100000010) && ({row_reg, col_reg}<18'b010010101100000100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010010101100000100)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b010010101100000101) && ({row_reg, col_reg}<18'b010010101100001000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010010101100001000) && ({row_reg, col_reg}<18'b010010101100001011)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b010010101100001011) && ({row_reg, col_reg}<18'b010010110000000010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010010110000000010) && ({row_reg, col_reg}<18'b010010110000000100)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}>=18'b010010110000000100) && ({row_reg, col_reg}<18'b010010110000000110)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==18'b010010110000000110)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}==18'b010010110000000111)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}>=18'b010010110000001000) && ({row_reg, col_reg}<18'b010010110000001010)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}>=18'b010010110000001010) && ({row_reg, col_reg}<18'b010010110000001101)) color_data = 12'b011011001101;
		if(({row_reg, col_reg}==18'b010010110000001101)) color_data = 12'b011111001110;
		if(({row_reg, col_reg}==18'b010010110000001110)) color_data = 12'b011011001110;
		if(({row_reg, col_reg}==18'b010010110000001111)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}>=18'b010010110000010000) && ({row_reg, col_reg}<18'b010010110000010010)) color_data = 12'b011110111110;
		if(({row_reg, col_reg}>=18'b010010110000010010) && ({row_reg, col_reg}<18'b010010110000010100)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}==18'b010010110000010100)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}==18'b010010110000010101)) color_data = 12'b010110101101;
		if(({row_reg, col_reg}==18'b010010110000010110)) color_data = 12'b011111011110;
		if(({row_reg, col_reg}>=18'b010010110000010111) && ({row_reg, col_reg}<18'b010010110000011010)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010010110000011010) && ({row_reg, col_reg}<18'b010010110000011100)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010010110000011100)) color_data = 12'b100011101110;
		if(({row_reg, col_reg}>=18'b010010110000011101) && ({row_reg, col_reg}<18'b010010110000100000)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010010110000100000)) color_data = 12'b010110101101;
		if(({row_reg, col_reg}>=18'b010010110000100001) && ({row_reg, col_reg}<18'b010010110000100011)) color_data = 12'b001110011100;
		if(({row_reg, col_reg}==18'b010010110000100011)) color_data = 12'b010010011011;
		if(({row_reg, col_reg}==18'b010010110000100100)) color_data = 12'b010110001010;
		if(({row_reg, col_reg}==18'b010010110000100101)) color_data = 12'b010101100111;
		if(({row_reg, col_reg}==18'b010010110000100110)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}==18'b010010110000100111)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010010110000101000) && ({row_reg, col_reg}<18'b010010110000101010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010010110000101010)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010010110000101011) && ({row_reg, col_reg}<18'b010010110000110010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010010110000110010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010010110000110011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010110000110100)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b010010110000110101) && ({row_reg, col_reg}<18'b010010110000111000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010110000111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010010110000111001)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b010010110000111010) && ({row_reg, col_reg}<18'b010010110000111100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010010110000111100)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}>=18'b010010110000111101) && ({row_reg, col_reg}<18'b010010110001000000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010010110001000000)) color_data = 12'b110010101011;
		if(({row_reg, col_reg}==18'b010010110001000001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010010110001000010) && ({row_reg, col_reg}<18'b010010110001000101)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010010110001000101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010010110001000110)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==18'b010010110001000111)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b010010110001001000) && ({row_reg, col_reg}<18'b010010110001001010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010010110001001010)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b010010110001001011) && ({row_reg, col_reg}<18'b010010110001001110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010110001001110)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==18'b010010110001001111)) color_data = 12'b011110011010;
		if(({row_reg, col_reg}>=18'b010010110001010000) && ({row_reg, col_reg}<18'b010010110001010100)) color_data = 12'b100011011111;
		if(({row_reg, col_reg}==18'b010010110001010100)) color_data = 12'b010110101110;
		if(({row_reg, col_reg}==18'b010010110001010101)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010010110001010110)) color_data = 12'b001010001110;
		if(({row_reg, col_reg}==18'b010010110001010111)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b010010110001011000)) color_data = 12'b001010001101;
		if(({row_reg, col_reg}==18'b010010110001011001)) color_data = 12'b011010111111;
		if(({row_reg, col_reg}>=18'b010010110001011010) && ({row_reg, col_reg}<18'b010010110001011101)) color_data = 12'b100011011111;
		if(({row_reg, col_reg}==18'b010010110001011101)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}==18'b010010110001011110)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010010110001011111)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}>=18'b010010110001100000) && ({row_reg, col_reg}<18'b010010110001100010)) color_data = 12'b100011011111;
		if(({row_reg, col_reg}==18'b010010110001100010)) color_data = 12'b011111001110;
		if(({row_reg, col_reg}==18'b010010110001100011)) color_data = 12'b010010001010;
		if(({row_reg, col_reg}==18'b010010110001100100)) color_data = 12'b010001111001;
		if(({row_reg, col_reg}==18'b010010110001100101)) color_data = 12'b010101111000;
		if(({row_reg, col_reg}==18'b010010110001100110)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==18'b010010110001100111)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}==18'b010010110001101000)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010010110001101001) && ({row_reg, col_reg}<18'b010010110001101100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010010110001101100)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}>=18'b010010110001101101) && ({row_reg, col_reg}<18'b010010110001110011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010010110001110011)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010010110001110100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010010110001110101)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010010110001110110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010010110001110111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010010110001111000) && ({row_reg, col_reg}<18'b010010110001111100)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==18'b010010110001111100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010010110001111101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010010110001111110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010010110001111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010010110010000000) && ({row_reg, col_reg}<18'b010010110010000100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010010110010000100)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==18'b010010110010000101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010010110010000110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010010110010000111)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==18'b010010110010001000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010010110010001001)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010010110010001010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010010110010001011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b010010110010001100) && ({row_reg, col_reg}<18'b010010110010001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010010110010001111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010010110010010000)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010010110010010001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010010110010010010)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b010010110010010011) && ({row_reg, col_reg}<18'b010010110010010111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010110010010111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010010110010011000) && ({row_reg, col_reg}<18'b010010110010011011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010010110010011011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010110010011100)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b010010110010011101) && ({row_reg, col_reg}<18'b010010110010011111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010010110010011111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010010110010100000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010010110010100001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010010110010100010)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010010110010100011) && ({row_reg, col_reg}<18'b010010110010100101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010010110010100101)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b010010110010100110) && ({row_reg, col_reg}<18'b010010110010110000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010110010110000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010010110010110001) && ({row_reg, col_reg}<18'b010010110010110100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010010110010110100) && ({row_reg, col_reg}<18'b010010110010111000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010010110010111000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010010110010111001)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}>=18'b010010110010111010) && ({row_reg, col_reg}<18'b010010110010111100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010010110010111100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010010110010111101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010010110010111110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010010110010111111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010110011000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010010110011000001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010010110011000010) && ({row_reg, col_reg}<18'b010010110011000110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010010110011000110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010010110011000111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010010110011001000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010010110011001001) && ({row_reg, col_reg}<18'b010010110011100011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010010110011100011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010010110011100100) && ({row_reg, col_reg}<18'b010010110011101000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010010110011101000)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010010110011101001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010010110011101010)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b010010110011101011) && ({row_reg, col_reg}<18'b010010110011110000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010010110011110000)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b010010110011110001) && ({row_reg, col_reg}<18'b010010110011110011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010010110011110011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010010110011110100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010010110011110101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010010110011110110)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010010110011110111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010010110011111000) && ({row_reg, col_reg}<18'b010010110011111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010010110011111010)) color_data = 12'b011110001000;
		if(({row_reg, col_reg}==18'b010010110011111011)) color_data = 12'b100010011010;
		if(({row_reg, col_reg}==18'b010010110011111100)) color_data = 12'b100010011011;
		if(({row_reg, col_reg}>=18'b010010110011111101) && ({row_reg, col_reg}<18'b010010110100000000)) color_data = 12'b011110011100;
		if(({row_reg, col_reg}>=18'b010010110100000000) && ({row_reg, col_reg}<18'b010010110100000010)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b010010110100000010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010010110100000011) && ({row_reg, col_reg}<18'b010010110100001000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010010110100001000) && ({row_reg, col_reg}<18'b010010110100001011)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b010010110100001011) && ({row_reg, col_reg}<18'b010010111000000000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010010111000000000)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}==18'b010010111000000001)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}==18'b010010111000000010)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==18'b010010111000000011)) color_data = 12'b100011011111;
		if(({row_reg, col_reg}==18'b010010111000000100)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b010010111000000101)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010010111000000110)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}>=18'b010010111000000111) && ({row_reg, col_reg}<18'b010010111000001001)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010010111000001001)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010010111000001010)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010010111000001011)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010010111000001100) && ({row_reg, col_reg}<18'b010010111000001110)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}>=18'b010010111000001110) && ({row_reg, col_reg}<18'b010010111000010000)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b010010111000010000)) color_data = 12'b101011101111;
		if(({row_reg, col_reg}==18'b010010111000010001)) color_data = 12'b100111011111;
		if(({row_reg, col_reg}==18'b010010111000010010)) color_data = 12'b011110111110;
		if(({row_reg, col_reg}>=18'b010010111000010011) && ({row_reg, col_reg}<18'b010010111000010101)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}==18'b010010111000010101)) color_data = 12'b010110101101;
		if(({row_reg, col_reg}==18'b010010111000010110)) color_data = 12'b011111011110;
		if(({row_reg, col_reg}>=18'b010010111000010111) && ({row_reg, col_reg}<18'b010010111000011011)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010010111000011011)) color_data = 12'b011011011101;
		if(({row_reg, col_reg}>=18'b010010111000011100) && ({row_reg, col_reg}<18'b010010111000011110)) color_data = 12'b011011001101;
		if(({row_reg, col_reg}==18'b010010111000011110)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}==18'b010010111000011111)) color_data = 12'b011011001110;
		if(({row_reg, col_reg}==18'b010010111000100000)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}>=18'b010010111000100001) && ({row_reg, col_reg}<18'b010010111000100011)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010010111000100011)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b010010111000100100)) color_data = 12'b100111001101;
		if(({row_reg, col_reg}==18'b010010111000100101)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==18'b010010111000100110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010010111000100111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010010111000101000) && ({row_reg, col_reg}<18'b010010111000101010)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==18'b010010111000101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010010111000101011) && ({row_reg, col_reg}<18'b010010111000110011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010010111000110011) && ({row_reg, col_reg}<18'b010010111000110111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010111000110111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010010111000111000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010010111000111001) && ({row_reg, col_reg}<18'b010010111000111011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010010111000111011)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010010111000111100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010010111000111101) && ({row_reg, col_reg}<18'b010010111001000001)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010010111001000001)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010010111001000010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010010111001000011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010111001000100)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010010111001000101)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010010111001000110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010010111001000111) && ({row_reg, col_reg}<18'b010010111001001010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010010111001001010)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010010111001001011)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==18'b010010111001001100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010111001001101)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}==18'b010010111001001110)) color_data = 12'b011001111000;
		if(({row_reg, col_reg}==18'b010010111001001111)) color_data = 12'b011010001000;
		if(({row_reg, col_reg}==18'b010010111001010000)) color_data = 12'b010010011011;
		if(({row_reg, col_reg}==18'b010010111001010001)) color_data = 12'b010010001011;
		if(({row_reg, col_reg}>=18'b010010111001010010) && ({row_reg, col_reg}<18'b010010111001010100)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b010010111001010100)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b010010111001010101)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010010111001010110) && ({row_reg, col_reg}<18'b010010111001011000)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b010010111001011000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010010111001011001)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}>=18'b010010111001011010) && ({row_reg, col_reg}<18'b010010111001011100)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b010010111001011100)) color_data = 12'b001110001011;
		if(({row_reg, col_reg}>=18'b010010111001011101) && ({row_reg, col_reg}<18'b010010111001011111)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b010010111001011111)) color_data = 12'b001110001011;
		if(({row_reg, col_reg}>=18'b010010111001100000) && ({row_reg, col_reg}<18'b010010111001100010)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}>=18'b010010111001100010) && ({row_reg, col_reg}<18'b010010111001100100)) color_data = 12'b001101111011;
		if(({row_reg, col_reg}==18'b010010111001100100)) color_data = 12'b010001111011;
		if(({row_reg, col_reg}==18'b010010111001100101)) color_data = 12'b010001111001;
		if(({row_reg, col_reg}==18'b010010111001100110)) color_data = 12'b010101111001;
		if(({row_reg, col_reg}==18'b010010111001100111)) color_data = 12'b011001111000;
		if(({row_reg, col_reg}==18'b010010111001101000)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}==18'b010010111001101001)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010010111001101010) && ({row_reg, col_reg}<18'b010010111001101111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010010111001101111)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010010111001110000) && ({row_reg, col_reg}<18'b010010111001110011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010010111001110011)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010010111001110100)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==18'b010010111001110101)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010010111001110110) && ({row_reg, col_reg}<18'b010010111010000000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010010111010000000) && ({row_reg, col_reg}<18'b010010111010000011)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}==18'b010010111010000011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010010111010000100) && ({row_reg, col_reg}<18'b010010111010000111)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010010111010000111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010111010001000)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b010010111010001001) && ({row_reg, col_reg}<18'b010010111010001011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010010111010001011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010010111010001100) && ({row_reg, col_reg}<18'b010010111010010000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010010111010010000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010010111010010001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010010111010010010)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b010010111010010011) && ({row_reg, col_reg}<18'b010010111010010111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010010111010010111) && ({row_reg, col_reg}<18'b010010111010011100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010010111010011100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010111010011101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010010111010011110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010111010011111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010010111010100000) && ({row_reg, col_reg}<18'b010010111010100010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010111010100010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010010111010100011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010111010100100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010010111010100101)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b010010111010100110) && ({row_reg, col_reg}<18'b010010111010101111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010111010101111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010010111010110000) && ({row_reg, col_reg}<18'b010010111010110011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010010111010110011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010010111010110100) && ({row_reg, col_reg}<18'b010010111010111000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010010111010111000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010010111010111001) && ({row_reg, col_reg}<18'b010010111010111101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010010111010111101)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b010010111010111110) && ({row_reg, col_reg}<18'b010010111011000001)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010010111011000001)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010010111011000010) && ({row_reg, col_reg}<18'b010010111011000110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010010111011000110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010010111011000111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010010111011001000) && ({row_reg, col_reg}<18'b010010111011001010)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010010111011001010) && ({row_reg, col_reg}<18'b010010111011001100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010010111011001100) && ({row_reg, col_reg}<18'b010010111011100111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010010111011100111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010010111011101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010010111011101001) && ({row_reg, col_reg}<18'b010010111011101011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010010111011101011) && ({row_reg, col_reg}<18'b010010111011101110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010010111011101110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010010111011101111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010010111011110000)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010010111011110001)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010010111011110010) && ({row_reg, col_reg}<18'b010010111011111000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010010111011111000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010010111011111001)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010010111011111010)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}>=18'b010010111011111011) && ({row_reg, col_reg}<18'b010010111011111101)) color_data = 12'b011001111000;
		if(({row_reg, col_reg}==18'b010010111011111101)) color_data = 12'b011001111001;
		if(({row_reg, col_reg}==18'b010010111011111110)) color_data = 12'b010101111001;
		if(({row_reg, col_reg}==18'b010010111011111111)) color_data = 12'b011010001010;
		if(({row_reg, col_reg}==18'b010010111100000000)) color_data = 12'b011110011100;
		if(({row_reg, col_reg}>=18'b010010111100000001) && ({row_reg, col_reg}<18'b010010111100000011)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b010010111100000011) && ({row_reg, col_reg}<18'b010010111100001000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010010111100001000) && ({row_reg, col_reg}<18'b010010111100001011)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b010010111100001011) && ({row_reg, col_reg}<18'b010011000000000000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010011000000000000)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}>=18'b010011000000000001) && ({row_reg, col_reg}<18'b010011000000000011)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}==18'b010011000000000011)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}==18'b010011000000000100)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b010011000000000101)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010011000000000110) && ({row_reg, col_reg}<18'b010011000000001011)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010011000000001011) && ({row_reg, col_reg}<18'b010011000000010000)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010011000000010000)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}==18'b010011000000010001)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b010011000000010010)) color_data = 12'b011110111101;
		if(({row_reg, col_reg}==18'b010011000000010011)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}==18'b010011000000010100)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}==18'b010011000000010101)) color_data = 12'b010110101101;
		if(({row_reg, col_reg}==18'b010011000000010110)) color_data = 12'b011111001110;
		if(({row_reg, col_reg}>=18'b010011000000010111) && ({row_reg, col_reg}<18'b010011000000011001)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}>=18'b010011000000011001) && ({row_reg, col_reg}<18'b010011000000011011)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010011000000011011)) color_data = 12'b011011001101;
		if(({row_reg, col_reg}>=18'b010011000000011100) && ({row_reg, col_reg}<18'b010011000000100000)) color_data = 12'b010110111101;
		if(({row_reg, col_reg}==18'b010011000000100000)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}>=18'b010011000000100001) && ({row_reg, col_reg}<18'b010011000000100011)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010011000000100011)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}==18'b010011000000100100)) color_data = 12'b101011011101;
		if(({row_reg, col_reg}==18'b010011000000100101)) color_data = 12'b010101110111;
		if(({row_reg, col_reg}==18'b010011000000100110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010011000000100111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011000000101000)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010011000000101001) && ({row_reg, col_reg}<18'b010011000000101011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010011000000101011) && ({row_reg, col_reg}<18'b010011000000101111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011000000101111)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010011000000110000) && ({row_reg, col_reg}<18'b010011000000110011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011000000110011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010011000000110100) && ({row_reg, col_reg}<18'b010011000000110110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010011000000110110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010011000000110111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010011000000111000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010011000000111001)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==18'b010011000000111010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010011000000111011)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}>=18'b010011000000111100) && ({row_reg, col_reg}<18'b010011000001000001)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010011000001000001)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b010011000001000010) && ({row_reg, col_reg}<18'b010011000001000100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010011000001000100) && ({row_reg, col_reg}<18'b010011000001000110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010011000001000110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010011000001000111)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==18'b010011000001001000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010011000001001001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==18'b010011000001001010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010011000001001011)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010011000001001100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010011000001001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010011000001001110)) color_data = 12'b011001111000;
		if(({row_reg, col_reg}==18'b010011000001001111)) color_data = 12'b011010001001;
		if(({row_reg, col_reg}==18'b010011000001010000)) color_data = 12'b001001111010;
		if(({row_reg, col_reg}==18'b010011000001010001)) color_data = 12'b001101111011;
		if(({row_reg, col_reg}==18'b010011000001010010)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}>=18'b010011000001010011) && ({row_reg, col_reg}<18'b010011000001010101)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010011000001010101)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b010011000001010110) && ({row_reg, col_reg}<18'b010011000001011000)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b010011000001011000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010011000001011001)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010011000001011010)) color_data = 12'b001001101011;
		if(({row_reg, col_reg}>=18'b010011000001011011) && ({row_reg, col_reg}<18'b010011000001100000)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}>=18'b010011000001100000) && ({row_reg, col_reg}<18'b010011000001100010)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010011000001100010)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b010011000001100011) && ({row_reg, col_reg}<18'b010011000001100101)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010011000001100101)) color_data = 12'b010001111011;
		if(({row_reg, col_reg}==18'b010011000001100110)) color_data = 12'b010001111010;
		if(({row_reg, col_reg}==18'b010011000001100111)) color_data = 12'b010101111001;
		if(({row_reg, col_reg}==18'b010011000001101000)) color_data = 12'b011001101000;
		if(({row_reg, col_reg}==18'b010011000001101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010011000001101010)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}>=18'b010011000001101011) && ({row_reg, col_reg}<18'b010011000001101101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011000001101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010011000001101110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011000001101111)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010011000001110000) && ({row_reg, col_reg}<18'b010011000001110010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011000001110010)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010011000001110011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011000001110100)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}>=18'b010011000001110101) && ({row_reg, col_reg}<18'b010011000001111001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010011000001111001)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}>=18'b010011000001111010) && ({row_reg, col_reg}<18'b010011000001111110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010011000001111110)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}>=18'b010011000001111111) && ({row_reg, col_reg}<18'b010011000010000100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010011000010000100) && ({row_reg, col_reg}<18'b010011000010000110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010011000010000110) && ({row_reg, col_reg}<18'b010011000010001001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010011000010001001) && ({row_reg, col_reg}<18'b010011000010010010)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010011000010010010)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b010011000010010011) && ({row_reg, col_reg}<18'b010011000010010111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010011000010010111) && ({row_reg, col_reg}<18'b010011000010011100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010011000010011100) && ({row_reg, col_reg}<18'b010011000010100011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010011000010100011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010011000010100100) && ({row_reg, col_reg}<18'b010011000010100111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010011000010100111)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b010011000010101000) && ({row_reg, col_reg}<18'b010011000010101110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010011000010101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010011000010101111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011000010110000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010011000010110001) && ({row_reg, col_reg}<18'b010011000010110011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011000010110011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010011000010110100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010011000010110101) && ({row_reg, col_reg}<18'b010011000010111000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010011000010111000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010011000010111001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010011000010111010) && ({row_reg, col_reg}<18'b010011000010111101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010011000010111101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010011000010111110) && ({row_reg, col_reg}<18'b010011000011000110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011000011000110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010011000011000111) && ({row_reg, col_reg}<18'b010011000011001011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010011000011001011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010011000011001100) && ({row_reg, col_reg}<18'b010011000011100111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010011000011100111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010011000011101000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010011000011101001) && ({row_reg, col_reg}<18'b010011000011101011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010011000011101011) && ({row_reg, col_reg}<18'b010011000011110011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010011000011110011) && ({row_reg, col_reg}<18'b010011000011110101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010011000011110101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010011000011110110) && ({row_reg, col_reg}<18'b010011000011111000)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010011000011111000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010011000011111001)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010011000011111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010011000011111011)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}==18'b010011000011111100)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==18'b010011000011111101)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}==18'b010011000011111110)) color_data = 12'b010101101000;
		if(({row_reg, col_reg}==18'b010011000011111111)) color_data = 12'b011001111001;
		if(({row_reg, col_reg}==18'b010011000100000000)) color_data = 12'b011110011100;
		if(({row_reg, col_reg}>=18'b010011000100000001) && ({row_reg, col_reg}<18'b010011000100000011)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b010011000100000011)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010011000100000100) && ({row_reg, col_reg}<18'b010011000100000111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010011000100000111) && ({row_reg, col_reg}<18'b010011000100001011)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b010011000100001011) && ({row_reg, col_reg}<18'b010011001000000000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010011001000000000) && ({row_reg, col_reg}<18'b010011001000000011)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}==18'b010011001000000011)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}==18'b010011001000000100)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}>=18'b010011001000000101) && ({row_reg, col_reg}<18'b010011001000000111)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010011001000000111) && ({row_reg, col_reg}<18'b010011001000001100)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010011001000001100) && ({row_reg, col_reg}<18'b010011001000010000)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010011001000010000)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}==18'b010011001000010001)) color_data = 12'b100011011111;
		if(({row_reg, col_reg}==18'b010011001000010010)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}>=18'b010011001000010011) && ({row_reg, col_reg}<18'b010011001000010101)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==18'b010011001000010101)) color_data = 12'b010110101101;
		if(({row_reg, col_reg}==18'b010011001000010110)) color_data = 12'b011111001111;
		if(({row_reg, col_reg}>=18'b010011001000010111) && ({row_reg, col_reg}<18'b010011001000011001)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}>=18'b010011001000011001) && ({row_reg, col_reg}<18'b010011001000011011)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010011001000011011)) color_data = 12'b011111011110;
		if(({row_reg, col_reg}>=18'b010011001000011100) && ({row_reg, col_reg}<18'b010011001000011111)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}==18'b010011001000011111)) color_data = 12'b010110111101;
		if(({row_reg, col_reg}>=18'b010011001000100000) && ({row_reg, col_reg}<18'b010011001000100011)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010011001000100011)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b010011001000100100)) color_data = 12'b101011011101;
		if(({row_reg, col_reg}==18'b010011001000100101)) color_data = 12'b010101110110;
		if(({row_reg, col_reg}==18'b010011001000100110)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}==18'b010011001000100111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010011001000101000)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010011001000101001) && ({row_reg, col_reg}<18'b010011001000101011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010011001000101011) && ({row_reg, col_reg}<18'b010011001000101111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011001000101111)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010011001000110000) && ({row_reg, col_reg}<18'b010011001000110011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011001000110011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010011001000110100) && ({row_reg, col_reg}<18'b010011001000110110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010011001000110110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010011001000110111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010011001000111000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010011001000111001)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010011001000111010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010011001000111011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010011001000111100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010011001000111101) && ({row_reg, col_reg}<18'b010011001001000000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010011001001000000)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==18'b010011001001000001)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==18'b010011001001000010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010011001001000011) && ({row_reg, col_reg}<18'b010011001001000101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010011001001000101)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010011001001000110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010011001001000111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==18'b010011001001001000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010011001001001001)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010011001001001010)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b010011001001001011) && ({row_reg, col_reg}<18'b010011001001001101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010011001001001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010011001001001110)) color_data = 12'b011110001001;
		if(({row_reg, col_reg}==18'b010011001001001111)) color_data = 12'b011010001010;
		if(({row_reg, col_reg}>=18'b010011001001010000) && ({row_reg, col_reg}<18'b010011001001010010)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b010011001001010010)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b010011001001010011)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b010011001001010100) && ({row_reg, col_reg}<18'b010011001001010111)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010011001001010111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010011001001011000)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}==18'b010011001001011001)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b010011001001011010)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010011001001011011)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b010011001001011100)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}>=18'b010011001001011101) && ({row_reg, col_reg}<18'b010011001001011111)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b010011001001011111)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010011001001100000)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010011001001100001)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}>=18'b010011001001100010) && ({row_reg, col_reg}<18'b010011001001100100)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010011001001100100) && ({row_reg, col_reg}<18'b010011001001100110)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010011001001100110)) color_data = 12'b010001111100;
		if(({row_reg, col_reg}==18'b010011001001100111)) color_data = 12'b010001111011;
		if(({row_reg, col_reg}==18'b010011001001101000)) color_data = 12'b010101111001;
		if(({row_reg, col_reg}>=18'b010011001001101001) && ({row_reg, col_reg}<18'b010011001001101011)) color_data = 12'b011001111000;
		if(({row_reg, col_reg}==18'b010011001001101011)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}>=18'b010011001001101100) && ({row_reg, col_reg}<18'b010011001001101110)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}==18'b010011001001101110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010011001001101111) && ({row_reg, col_reg}<18'b010011001001110100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010011001001110100) && ({row_reg, col_reg}<18'b010011001001110111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010011001001110111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010011001001111000) && ({row_reg, col_reg}<18'b010011001001111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010011001001111010)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010011001001111011) && ({row_reg, col_reg}<18'b010011001001111101)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010011001001111101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011001001111110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010011001001111111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010011001010000000)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==18'b010011001010000001)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}>=18'b010011001010000010) && ({row_reg, col_reg}<18'b010011001010000100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010011001010000100) && ({row_reg, col_reg}<18'b010011001010000110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010011001010000110) && ({row_reg, col_reg}<18'b010011001010001000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010011001010001000)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010011001010001001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010011001010001010)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b010011001010001011) && ({row_reg, col_reg}<18'b010011001010010000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010011001010010000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010011001010010001)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010011001010010010)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b010011001010010011) && ({row_reg, col_reg}<18'b010011001010010111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010011001010010111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010011001010011000) && ({row_reg, col_reg}<18'b010011001010011011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011001010011011)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010011001010011100) && ({row_reg, col_reg}<18'b010011001010101110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010011001010101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010011001010101111) && ({row_reg, col_reg}<18'b010011001010110011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011001010110011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010011001010110100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010011001010110101) && ({row_reg, col_reg}<18'b010011001010111000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010011001010111000)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010011001010111001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010011001010111010) && ({row_reg, col_reg}<18'b010011001010111101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010011001010111101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010011001010111110) && ({row_reg, col_reg}<18'b010011001011000110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011001011000110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010011001011000111) && ({row_reg, col_reg}<18'b010011001011001011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010011001011001011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010011001011001100) && ({row_reg, col_reg}<18'b010011001011101000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010011001011101000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010011001011101001) && ({row_reg, col_reg}<18'b010011001011110110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011001011110110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010011001011110111) && ({row_reg, col_reg}<18'b010011001011111011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010011001011111011) && ({row_reg, col_reg}<18'b010011001011111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010011001011111101)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}==18'b010011001011111110)) color_data = 12'b010101100111;
		if(({row_reg, col_reg}==18'b010011001011111111)) color_data = 12'b011001111001;
		if(({row_reg, col_reg}==18'b010011001100000000)) color_data = 12'b011110011100;
		if(({row_reg, col_reg}==18'b010011001100000001)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}==18'b010011001100000010)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b010011001100000011) && ({row_reg, col_reg}<18'b010011001100000101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010011001100000101) && ({row_reg, col_reg}<18'b010011001100001000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010011001100001000) && ({row_reg, col_reg}<18'b010011001100001011)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b010011001100001011) && ({row_reg, col_reg}<18'b010011010000000010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010011010000000010)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}==18'b010011010000000011)) color_data = 12'b100011011111;
		if(({row_reg, col_reg}==18'b010011010000000100)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}>=18'b010011010000000101) && ({row_reg, col_reg}<18'b010011010000001000)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010011010000001000) && ({row_reg, col_reg}<18'b010011010000001011)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010011010000001011) && ({row_reg, col_reg}<18'b010011010000010000)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010011010000010000)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}==18'b010011010000010001)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b010011010000010010)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}>=18'b010011010000010011) && ({row_reg, col_reg}<18'b010011010000010101)) color_data = 12'b011010111111;
		if(({row_reg, col_reg}==18'b010011010000010101)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==18'b010011010000010110)) color_data = 12'b011111001111;
		if(({row_reg, col_reg}>=18'b010011010000010111) && ({row_reg, col_reg}<18'b010011010000011001)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}>=18'b010011010000011001) && ({row_reg, col_reg}<18'b010011010000011011)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010011010000011011)) color_data = 12'b011011001110;
		if(({row_reg, col_reg}==18'b010011010000011100)) color_data = 12'b010110111101;
		if(({row_reg, col_reg}==18'b010011010000011101)) color_data = 12'b010110101100;
		if(({row_reg, col_reg}==18'b010011010000011110)) color_data = 12'b010110111101;
		if(({row_reg, col_reg}==18'b010011010000011111)) color_data = 12'b010110111100;
		if(({row_reg, col_reg}==18'b010011010000100000)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b010011010000100001)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010011010000100010) && ({row_reg, col_reg}<18'b010011010000100100)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}==18'b010011010000100100)) color_data = 12'b101011101110;
		if(({row_reg, col_reg}==18'b010011010000100101)) color_data = 12'b010101110110;
		if(({row_reg, col_reg}==18'b010011010000100110)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}>=18'b010011010000100111) && ({row_reg, col_reg}<18'b010011010000101001)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011010000101001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010011010000101010)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010011010000101011) && ({row_reg, col_reg}<18'b010011010000101111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011010000101111)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010011010000110000) && ({row_reg, col_reg}<18'b010011010000110011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011010000110011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010011010000110100) && ({row_reg, col_reg}<18'b010011010000110111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010011010000110111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010011010000111000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010011010000111001)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==18'b010011010000111010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010011010000111011)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=18'b010011010000111100) && ({row_reg, col_reg}<18'b010011010001000000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010011010001000000)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==18'b010011010001000001)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}>=18'b010011010001000010) && ({row_reg, col_reg}<18'b010011010001000101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010011010001000101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010011010001000110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010011010001000111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=18'b010011010001001000) && ({row_reg, col_reg}<18'b010011010001001011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010011010001001011)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==18'b010011010001001100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010011010001001101)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==18'b010011010001001110)) color_data = 12'b011001111001;
		if(({row_reg, col_reg}==18'b010011010001001111)) color_data = 12'b011010001010;
		if(({row_reg, col_reg}==18'b010011010001010000)) color_data = 12'b001001101100;
		if(({row_reg, col_reg}==18'b010011010001010001)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010011010001010010)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010011010001010011) && ({row_reg, col_reg}<18'b010011010001010101)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}>=18'b010011010001010101) && ({row_reg, col_reg}<18'b010011010001010111)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b010011010001010111) && ({row_reg, col_reg}<18'b010011010001011001)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010011010001011001) && ({row_reg, col_reg}<18'b010011010001011011)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010011010001011011)) color_data = 12'b001101111011;
		if(({row_reg, col_reg}==18'b010011010001011100)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}>=18'b010011010001011101) && ({row_reg, col_reg}<18'b010011010001011111)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010011010001011111)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}>=18'b010011010001100000) && ({row_reg, col_reg}<18'b010011010001100011)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010011010001100011)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010011010001100100) && ({row_reg, col_reg}<18'b010011010001100111)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010011010001100111)) color_data = 12'b010001111100;
		if(({row_reg, col_reg}==18'b010011010001101000)) color_data = 12'b010001111011;
		if(({row_reg, col_reg}==18'b010011010001101001)) color_data = 12'b010001111010;
		if(({row_reg, col_reg}==18'b010011010001101010)) color_data = 12'b010101111001;
		if(({row_reg, col_reg}==18'b010011010001101011)) color_data = 12'b010101101000;
		if(({row_reg, col_reg}==18'b010011010001101100)) color_data = 12'b011001101000;
		if(({row_reg, col_reg}==18'b010011010001101101)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==18'b010011010001101110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010011010001101111) && ({row_reg, col_reg}<18'b010011010001110010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010011010001110010) && ({row_reg, col_reg}<18'b010011010001110110)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}>=18'b010011010001110110) && ({row_reg, col_reg}<18'b010011010001111001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010011010001111001)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011010001111010)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==18'b010011010001111011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010011010001111100) && ({row_reg, col_reg}<18'b010011010001111110)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}>=18'b010011010001111110) && ({row_reg, col_reg}<18'b010011010010000000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011010010000000)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==18'b010011010010000001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010011010010000010) && ({row_reg, col_reg}<18'b010011010010000100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011010010000100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010011010010000101) && ({row_reg, col_reg}<18'b010011010010001001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010011010010001001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b010011010010001010) && ({row_reg, col_reg}<18'b010011010010010010)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010011010010010010)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b010011010010010011) && ({row_reg, col_reg}<18'b010011010010010111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010011010010010111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010011010010011000) && ({row_reg, col_reg}<18'b010011010010011011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011010010011011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010011010010011100) && ({row_reg, col_reg}<18'b010011010010101111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010011010010101111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010011010010110000) && ({row_reg, col_reg}<18'b010011010010110011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011010010110011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010011010010110100) && ({row_reg, col_reg}<18'b010011010010111000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010011010010111000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010011010010111001) && ({row_reg, col_reg}<18'b010011010010111011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010011010010111011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010011010010111100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010011010010111101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010011010010111110) && ({row_reg, col_reg}<18'b010011010011000110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011010011000110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010011010011000111) && ({row_reg, col_reg}<18'b010011010011001011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010011010011001011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010011010011001100) && ({row_reg, col_reg}<18'b010011010011100111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010011010011100111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010011010011101000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010011010011101001) && ({row_reg, col_reg}<18'b010011010011101100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011010011101100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010011010011101101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011010011101110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010011010011101111) && ({row_reg, col_reg}<18'b010011010011110110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011010011110110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010011010011110111) && ({row_reg, col_reg}<18'b010011010011111010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010011010011111010)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==18'b010011010011111011)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010011010011111100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011010011111101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010011010011111110)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}==18'b010011010011111111)) color_data = 12'b011001111000;
		if(({row_reg, col_reg}==18'b010011010100000000)) color_data = 12'b011110011100;
		if(({row_reg, col_reg}==18'b010011010100000001)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b010011010100000010) && ({row_reg, col_reg}<18'b010011010100000100)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b010011010100000100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010011010100000101) && ({row_reg, col_reg}<18'b010011010100000111)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b010011010100000111) && ({row_reg, col_reg}<18'b010011010100001011)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b010011010100001011) && ({row_reg, col_reg}<18'b010011011000000010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010011011000000010)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==18'b010011011000000011)) color_data = 12'b011111001110;
		if(({row_reg, col_reg}==18'b010011011000000100)) color_data = 12'b011111001111;
		if(({row_reg, col_reg}>=18'b010011011000000101) && ({row_reg, col_reg}<18'b010011011000001000)) color_data = 12'b011111001110;
		if(({row_reg, col_reg}>=18'b010011011000001000) && ({row_reg, col_reg}<18'b010011011000001101)) color_data = 12'b011111011110;
		if(({row_reg, col_reg}==18'b010011011000001101)) color_data = 12'b100011011110;
		if(({row_reg, col_reg}==18'b010011011000001110)) color_data = 12'b011111011110;
		if(({row_reg, col_reg}==18'b010011011000001111)) color_data = 12'b011111001110;
		if(({row_reg, col_reg}==18'b010011011000010000)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}==18'b010011011000010001)) color_data = 12'b011111001110;
		if(({row_reg, col_reg}==18'b010011011000010010)) color_data = 12'b010110011101;
		if(({row_reg, col_reg}>=18'b010011011000010011) && ({row_reg, col_reg}<18'b010011011000010110)) color_data = 12'b010010011101;
		if(({row_reg, col_reg}>=18'b010011011000010110) && ({row_reg, col_reg}<18'b010011011000011000)) color_data = 12'b010110101110;
		if(({row_reg, col_reg}==18'b010011011000011000)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}>=18'b010011011000011001) && ({row_reg, col_reg}<18'b010011011000011011)) color_data = 12'b010110111101;
		if(({row_reg, col_reg}==18'b010011011000011011)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}==18'b010011011000011100)) color_data = 12'b100011011111;
		if(({row_reg, col_reg}==18'b010011011000011101)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}==18'b010011011000011110)) color_data = 12'b100011011111;
		if(({row_reg, col_reg}==18'b010011011000011111)) color_data = 12'b011111011110;
		if(({row_reg, col_reg}>=18'b010011011000100000) && ({row_reg, col_reg}<18'b010011011000100010)) color_data = 12'b010110111101;
		if(({row_reg, col_reg}==18'b010011011000100010)) color_data = 12'b010110111110;
		if(({row_reg, col_reg}==18'b010011011000100011)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}==18'b010011011000100100)) color_data = 12'b011010011011;
		if(({row_reg, col_reg}==18'b010011011000100101)) color_data = 12'b011001111000;
		if(({row_reg, col_reg}==18'b010011011000100110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010011011000100111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011011000101000)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010011011000101001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010011011000101010)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010011011000101011) && ({row_reg, col_reg}<18'b010011011000101111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011011000101111)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010011011000110000) && ({row_reg, col_reg}<18'b010011011000110011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011011000110011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010011011000110100) && ({row_reg, col_reg}<18'b010011011000110111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010011011000110111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010011011000111000)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010011011000111001)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==18'b010011011000111010)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010011011000111011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b010011011000111100) && ({row_reg, col_reg}<18'b010011011000111110)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010011011000111110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010011011000111111)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010011011001000000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010011011001000001)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b010011011001000010) && ({row_reg, col_reg}<18'b010011011001000101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010011011001000101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010011011001000110) && ({row_reg, col_reg}<18'b010011011001001000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010011011001001000) && ({row_reg, col_reg}<18'b010011011001001011)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010011011001001011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010011011001001100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011011001001101)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==18'b010011011001001110)) color_data = 12'b011001111000;
		if(({row_reg, col_reg}==18'b010011011001001111)) color_data = 12'b010101111001;
		if(({row_reg, col_reg}==18'b010011011001010000)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b010011011001010001) && ({row_reg, col_reg}<18'b010011011001010011)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010011011001010011)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b010011011001010100)) color_data = 12'b001101111111;
		if(({row_reg, col_reg}==18'b010011011001010101)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b010011011001010110)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010011011001010111)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}==18'b010011011001011000)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010011011001011001)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b010011011001011010)) color_data = 12'b011110111111;
		if(({row_reg, col_reg}==18'b010011011001011011)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==18'b010011011001011100)) color_data = 12'b011011001111;
		if(({row_reg, col_reg}==18'b010011011001011101)) color_data = 12'b011011001110;
		if(({row_reg, col_reg}==18'b010011011001011110)) color_data = 12'b011011001111;
		if(({row_reg, col_reg}>=18'b010011011001011111) && ({row_reg, col_reg}<18'b010011011001100001)) color_data = 12'b010111001110;
		if(({row_reg, col_reg}==18'b010011011001100001)) color_data = 12'b011011001111;
		if(({row_reg, col_reg}==18'b010011011001100010)) color_data = 12'b010110111110;
		if(({row_reg, col_reg}==18'b010011011001100011)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010011011001100100)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010011011001100101)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b010011011001100110) && ({row_reg, col_reg}<18'b010011011001101000)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010011011001101000)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010011011001101001)) color_data = 12'b010001111011;
		if(({row_reg, col_reg}==18'b010011011001101010)) color_data = 12'b010001111010;
		if(({row_reg, col_reg}==18'b010011011001101011)) color_data = 12'b010101111001;
		if(({row_reg, col_reg}==18'b010011011001101100)) color_data = 12'b011110001010;
		if(({row_reg, col_reg}==18'b010011011001101101)) color_data = 12'b100010011010;
		if(({row_reg, col_reg}==18'b010011011001101110)) color_data = 12'b100110001001;
		if(({row_reg, col_reg}==18'b010011011001101111)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010011011001110000)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==18'b010011011001110001)) color_data = 12'b101010011000;
		if(({row_reg, col_reg}==18'b010011011001110010)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}>=18'b010011011001110011) && ({row_reg, col_reg}<18'b010011011001110110)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010011011001110110)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==18'b010011011001110111)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010011011001111000)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}>=18'b010011011001111001) && ({row_reg, col_reg}<18'b010011011001111011)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010011011001111011)) color_data = 12'b101010001000;
		if(({row_reg, col_reg}>=18'b010011011001111100) && ({row_reg, col_reg}<18'b010011011001111110)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==18'b010011011001111110)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010011011001111111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010011011010000000) && ({row_reg, col_reg}<18'b010011011010000100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011011010000100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010011011010000101) && ({row_reg, col_reg}<18'b010011011010001000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010011011010001000)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b010011011010001001) && ({row_reg, col_reg}<18'b010011011010001011)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010011011010001011) && ({row_reg, col_reg}<18'b010011011010001110)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b010011011010001110) && ({row_reg, col_reg}<18'b010011011010010010)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010011011010010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010011011010010011) && ({row_reg, col_reg}<18'b010011011010010110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010011011010010110) && ({row_reg, col_reg}<18'b010011011010011011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011011010011011)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010011011010011100) && ({row_reg, col_reg}<18'b010011011010101001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010011011010101001) && ({row_reg, col_reg}<18'b010011011010101011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010011011010101011)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010011011010101100) && ({row_reg, col_reg}<18'b010011011010101110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010011011010101110) && ({row_reg, col_reg}<18'b010011011010110011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011011010110011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010011011010110100) && ({row_reg, col_reg}<18'b010011011010110110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010011011010110110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010011011010110111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010011011010111000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010011011010111001) && ({row_reg, col_reg}<18'b010011011010111011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010011011010111011)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010011011010111100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010011011010111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010011011010111110) && ({row_reg, col_reg}<18'b010011011011000001)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011011011000001)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010011011011000010) && ({row_reg, col_reg}<18'b010011011011000110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011011011000110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010011011011000111) && ({row_reg, col_reg}<18'b010011011011001001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010011011011001001)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010011011011001010)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010011011011001011)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b010011011011001100) && ({row_reg, col_reg}<18'b010011011011001110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010011011011001110) && ({row_reg, col_reg}<18'b010011011011010000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010011011011010000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010011011011010001) && ({row_reg, col_reg}<18'b010011011011010011)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010011011011010011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b010011011011010100) && ({row_reg, col_reg}<18'b010011011011010110)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==18'b010011011011010110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010011011011010111)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==18'b010011011011011000)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010011011011011001)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}>=18'b010011011011011010) && ({row_reg, col_reg}<18'b010011011011011101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010011011011011101)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}>=18'b010011011011011110) && ({row_reg, col_reg}<18'b010011011011100000)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010011011011100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010011011011100001) && ({row_reg, col_reg}<18'b010011011011100111)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010011011011100111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010011011011101000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010011011011101001) && ({row_reg, col_reg}<18'b010011011011110110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011011011110110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010011011011110111) && ({row_reg, col_reg}<18'b010011011011111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010011011011111010)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}>=18'b010011011011111011) && ({row_reg, col_reg}<18'b010011011011111110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010011011011111110) && ({row_reg, col_reg}<18'b010011011100000000)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}==18'b010011011100000000)) color_data = 12'b011110011100;
		if(({row_reg, col_reg}==18'b010011011100000001)) color_data = 12'b011110011101;
		if(({row_reg, col_reg}>=18'b010011011100000010) && ({row_reg, col_reg}<18'b010011011100000100)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b010011011100000100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010011011100000101) && ({row_reg, col_reg}<18'b010011011100000111)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b010011011100000111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010011011100001000) && ({row_reg, col_reg}<18'b010011011100001011)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b010011011100001011) && ({row_reg, col_reg}<18'b010011100000000100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010011100000000100) && ({row_reg, col_reg}<18'b010011100000001001)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}==18'b010011100000001001)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}>=18'b010011100000001010) && ({row_reg, col_reg}<18'b010011100000001101)) color_data = 12'b010110101101;
		if(({row_reg, col_reg}==18'b010011100000001101)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}==18'b010011100000001110)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}==18'b010011100000001111)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}==18'b010011100000010000)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==18'b010011100000010001)) color_data = 12'b010110101101;
		if(({row_reg, col_reg}==18'b010011100000010010)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b010011100000010011)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}>=18'b010011100000010100) && ({row_reg, col_reg}<18'b010011100000010111)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b010011100000010111) && ({row_reg, col_reg}<18'b010011100000011001)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}>=18'b010011100000011001) && ({row_reg, col_reg}<18'b010011100000011011)) color_data = 12'b000101111010;
		if(({row_reg, col_reg}==18'b010011100000011011)) color_data = 12'b011011001110;
		if(({row_reg, col_reg}==18'b010011100000011100)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010011100000011101)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010011100000011110)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}==18'b010011100000011111)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010011100000100000)) color_data = 12'b010010011100;
		if(({row_reg, col_reg}==18'b010011100000100001)) color_data = 12'b001001111010;
		if(({row_reg, col_reg}==18'b010011100000100010)) color_data = 12'b000101101010;
		if(({row_reg, col_reg}==18'b010011100000100011)) color_data = 12'b001101111010;
		if(({row_reg, col_reg}==18'b010011100000100100)) color_data = 12'b010001111001;
		if(({row_reg, col_reg}==18'b010011100000100101)) color_data = 12'b010101110111;
		if(({row_reg, col_reg}==18'b010011100000100110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010011100000100111) && ({row_reg, col_reg}<18'b010011100000101001)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010011100000101001) && ({row_reg, col_reg}<18'b010011100000101100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010011100000101100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011100000101101)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010011100000101110) && ({row_reg, col_reg}<18'b010011100000110011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011100000110011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010011100000110100) && ({row_reg, col_reg}<18'b010011100000110110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010011100000110110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010011100000110111) && ({row_reg, col_reg}<18'b010011100000111001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010011100000111001)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b010011100000111010) && ({row_reg, col_reg}<18'b010011100000111100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010011100000111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010011100000111101) && ({row_reg, col_reg}<18'b010011100001000010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011100001000010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010011100001000011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011100001000100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010011100001000101) && ({row_reg, col_reg}<18'b010011100001001001)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011100001001001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010011100001001010) && ({row_reg, col_reg}<18'b010011100001001100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010011100001001100) && ({row_reg, col_reg}<18'b010011100001001110)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==18'b010011100001001110)) color_data = 12'b011001101000;
		if(({row_reg, col_reg}==18'b010011100001001111)) color_data = 12'b010101111001;
		if(({row_reg, col_reg}>=18'b010011100001010000) && ({row_reg, col_reg}<18'b010011100001010010)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010011100001010010)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010011100001010011)) color_data = 12'b001110001111;
		if(({row_reg, col_reg}==18'b010011100001010100)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}==18'b010011100001010101)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010011100001010110)) color_data = 12'b000101101100;
		if(({row_reg, col_reg}>=18'b010011100001010111) && ({row_reg, col_reg}<18'b010011100001011001)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010011100001011001)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}>=18'b010011100001011010) && ({row_reg, col_reg}<18'b010011100001011101)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010011100001011101) && ({row_reg, col_reg}<18'b010011100001100001)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010011100001100001)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010011100001100010)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}==18'b010011100001100011)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b010011100001100100)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010011100001100101)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b010011100001100110) && ({row_reg, col_reg}<18'b010011100001101000)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b010011100001101000) && ({row_reg, col_reg}<18'b010011100001101010)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010011100001101010)) color_data = 12'b010001111011;
		if(({row_reg, col_reg}==18'b010011100001101011)) color_data = 12'b010001111010;
		if(({row_reg, col_reg}==18'b010011100001101100)) color_data = 12'b100010011011;
		if(({row_reg, col_reg}==18'b010011100001101101)) color_data = 12'b101010111100;
		if(({row_reg, col_reg}==18'b010011100001101110)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b010011100001101111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010011100001110000) && ({row_reg, col_reg}<18'b010011100001110011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b010011100001110011) && ({row_reg, col_reg}<18'b010011100001110101)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}>=18'b010011100001110101) && ({row_reg, col_reg}<18'b010011100001110111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==18'b010011100001110111)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}>=18'b010011100001111000) && ({row_reg, col_reg}<18'b010011100001111010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010011100001111010)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==18'b010011100001111011)) color_data = 12'b110010111010;
		if(({row_reg, col_reg}==18'b010011100001111100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010011100001111101)) color_data = 12'b110010111010;
		if(({row_reg, col_reg}==18'b010011100001111110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010011100001111111)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b010011100010000000) && ({row_reg, col_reg}<18'b010011100010000100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011100010000100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010011100010000101) && ({row_reg, col_reg}<18'b010011100010000111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010011100010000111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010011100010001000) && ({row_reg, col_reg}<18'b010011100010001010)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b010011100010001010) && ({row_reg, col_reg}<18'b010011100010001100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010011100010001100)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010011100010001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010011100010001110) && ({row_reg, col_reg}<18'b010011100010010010)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010011100010010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010011100010010011) && ({row_reg, col_reg}<18'b010011100010011100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010011100010011100) && ({row_reg, col_reg}<18'b010011100010101010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010011100010101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010011100010101011) && ({row_reg, col_reg}<18'b010011100010110011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011100010110011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010011100010110100) && ({row_reg, col_reg}<18'b010011100010110110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010011100010110110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010011100010110111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010011100010111000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b010011100010111001) && ({row_reg, col_reg}<18'b010011100011000110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011100011000110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010011100011000111) && ({row_reg, col_reg}<18'b010011100011010000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010011100011010000)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b010011100011010001) && ({row_reg, col_reg}<18'b010011100011011110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010011100011011110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010011100011011111) && ({row_reg, col_reg}<18'b010011100011101010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011100011101010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010011100011101011) && ({row_reg, col_reg}<18'b010011100011110100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011100011110100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010011100011110101) && ({row_reg, col_reg}<18'b010011100011111011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011100011111011)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}>=18'b010011100011111100) && ({row_reg, col_reg}<18'b010011100011111110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011100011111110)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==18'b010011100011111111)) color_data = 12'b011001111000;
		if(({row_reg, col_reg}>=18'b010011100100000000) && ({row_reg, col_reg}<18'b010011100100000010)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}>=18'b010011100100000010) && ({row_reg, col_reg}<18'b010011100100000100)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010011100100000100) && ({row_reg, col_reg}<18'b010011100100000111)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b010011100100000111) && ({row_reg, col_reg}<18'b010011100100001001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010011100100001001) && ({row_reg, col_reg}<18'b010011100100001011)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b010011100100001011) && ({row_reg, col_reg}<18'b010011101000000101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010011101000000101) && ({row_reg, col_reg}<18'b010011101000001000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010011101000001000) && ({row_reg, col_reg}<18'b010011101000001100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010011101000001100)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}>=18'b010011101000001101) && ({row_reg, col_reg}<18'b010011101000010000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010011101000010000)) color_data = 12'b011010111111;
		if(({row_reg, col_reg}==18'b010011101000010001)) color_data = 12'b010110101110;
		if(({row_reg, col_reg}==18'b010011101000010010)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b010011101000010011)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b010011101000010100) && ({row_reg, col_reg}<18'b010011101000011000)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b010011101000011000)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b010011101000011001)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b010011101000011010)) color_data = 12'b000101111010;
		if(({row_reg, col_reg}==18'b010011101000011011)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}>=18'b010011101000011100) && ({row_reg, col_reg}<18'b010011101000011111)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010011101000011111)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010011101000100000)) color_data = 12'b010010101101;
		if(({row_reg, col_reg}==18'b010011101000100001)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b010011101000100010)) color_data = 12'b001110011100;
		if(({row_reg, col_reg}==18'b010011101000100011)) color_data = 12'b001101111011;
		if(({row_reg, col_reg}==18'b010011101000100100)) color_data = 12'b010110001011;
		if(({row_reg, col_reg}==18'b010011101000100101)) color_data = 12'b011001111000;
		if(({row_reg, col_reg}==18'b010011101000100110)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}==18'b010011101000100111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010011101000101000) && ({row_reg, col_reg}<18'b010011101000101011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010011101000101011) && ({row_reg, col_reg}<18'b010011101000110011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010011101000110011) && ({row_reg, col_reg}<18'b010011101000111100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010011101000111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010011101000111101) && ({row_reg, col_reg}<18'b010011101001000000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011101001000000)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010011101001000001) && ({row_reg, col_reg}<18'b010011101001001000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011101001001000)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010011101001001001) && ({row_reg, col_reg}<18'b010011101001001101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011101001001101)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==18'b010011101001001110)) color_data = 12'b011001101000;
		if(({row_reg, col_reg}==18'b010011101001001111)) color_data = 12'b010101111001;
		if(({row_reg, col_reg}>=18'b010011101001010000) && ({row_reg, col_reg}<18'b010011101001010011)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b010011101001010011) && ({row_reg, col_reg}<18'b010011101001010101)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010011101001010101)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b010011101001010110) && ({row_reg, col_reg}<18'b010011101001011000)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b010011101001011000)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b010011101001011001)) color_data = 12'b011111001111;
		if(({row_reg, col_reg}==18'b010011101001011010)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010011101001011011) && ({row_reg, col_reg}<18'b010011101001100001)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010011101001100001)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010011101001100010)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}==18'b010011101001100011)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}>=18'b010011101001100100) && ({row_reg, col_reg}<18'b010011101001100111)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010011101001100111)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b010011101001101000) && ({row_reg, col_reg}<18'b010011101001101010)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010011101001101010)) color_data = 12'b010001111010;
		if(({row_reg, col_reg}==18'b010011101001101011)) color_data = 12'b010001101001;
		if(({row_reg, col_reg}==18'b010011101001101100)) color_data = 12'b100010011011;
		if(({row_reg, col_reg}==18'b010011101001101101)) color_data = 12'b101010111100;
		if(({row_reg, col_reg}==18'b010011101001101110)) color_data = 12'b101010111011;
		if(({row_reg, col_reg}==18'b010011101001101111)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}>=18'b010011101001110000) && ({row_reg, col_reg}<18'b010011101001110010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010011101001110010) && ({row_reg, col_reg}<18'b010011101001111010)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}>=18'b010011101001111010) && ({row_reg, col_reg}<18'b010011101001111101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010011101001111101)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==18'b010011101001111110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010011101001111111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010011101010000000) && ({row_reg, col_reg}<18'b010011101010000010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010011101010000010) && ({row_reg, col_reg}<18'b010011101010000100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010011101010000100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010011101010000101) && ({row_reg, col_reg}<18'b010011101010001011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010011101010001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010011101010001100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010011101010001101)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010011101010001110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010011101010001111)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b010011101010010000) && ({row_reg, col_reg}<18'b010011101010010010)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010011101010010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010011101010010011) && ({row_reg, col_reg}<18'b010011101010011100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010011101010011100) && ({row_reg, col_reg}<18'b010011101010101010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010011101010101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010011101010101011) && ({row_reg, col_reg}<18'b010011101010110011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011101010110011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010011101010110100) && ({row_reg, col_reg}<18'b010011101010110110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010011101010110110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010011101010110111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010011101010111000)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010011101010111001)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011101010111010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010011101010111011) && ({row_reg, col_reg}<18'b010011101011000110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011101011000110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010011101011000111) && ({row_reg, col_reg}<18'b010011101011001001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010011101011001001)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b010011101011001010) && ({row_reg, col_reg}<18'b010011101011001100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010011101011001100)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b010011101011001101) && ({row_reg, col_reg}<18'b010011101011010000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010011101011010000)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b010011101011010001) && ({row_reg, col_reg}<18'b010011101011011110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010011101011011110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010011101011011111) && ({row_reg, col_reg}<18'b010011101011110011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010011101011110011) && ({row_reg, col_reg}<18'b010011101011110101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010011101011110101) && ({row_reg, col_reg}<18'b010011101011111011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010011101011111011) && ({row_reg, col_reg}<18'b010011101011111101)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==18'b010011101011111101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011101011111110)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==18'b010011101011111111)) color_data = 12'b011001111000;
		if(({row_reg, col_reg}==18'b010011101100000000)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}>=18'b010011101100000001) && ({row_reg, col_reg}<18'b010011101100000011)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b010011101100000011) && ({row_reg, col_reg}<18'b010011101100000101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010011101100000101) && ({row_reg, col_reg}<18'b010011101100001000)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b010011101100001000) && ({row_reg, col_reg}<18'b010011101100001100)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b010011101100001100) && ({row_reg, col_reg}<18'b010011110000000011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010011110000000011) && ({row_reg, col_reg}<18'b010011110000001100)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010011110000001100) && ({row_reg, col_reg}<18'b010011110000010000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010011110000010000)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b010011110000010001)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}>=18'b010011110000010010) && ({row_reg, col_reg}<18'b010011110000010100)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}>=18'b010011110000010100) && ({row_reg, col_reg}<18'b010011110000010111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010011110000010111)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010011110000011000)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010011110000011001)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b010011110000011010)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b010011110000011011)) color_data = 12'b011011001110;
		if(({row_reg, col_reg}>=18'b010011110000011100) && ({row_reg, col_reg}<18'b010011110000011111)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010011110000011111)) color_data = 12'b100011101110;
		if(({row_reg, col_reg}==18'b010011110000100000)) color_data = 12'b001110011100;
		if(({row_reg, col_reg}==18'b010011110000100001)) color_data = 12'b000101111010;
		if(({row_reg, col_reg}==18'b010011110000100010)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b010011110000100011)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b010011110000100100)) color_data = 12'b010001111010;
		if(({row_reg, col_reg}==18'b010011110000100101)) color_data = 12'b010101100111;
		if(({row_reg, col_reg}==18'b010011110000100110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010011110000100111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010011110000101000)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==18'b010011110000101001)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}>=18'b010011110000101010) && ({row_reg, col_reg}<18'b010011110000101100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010011110000101100) && ({row_reg, col_reg}<18'b010011110000101111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011110000101111)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010011110000110000) && ({row_reg, col_reg}<18'b010011110000110011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010011110000110011) && ({row_reg, col_reg}<18'b010011110000111011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010011110000111011)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010011110000111100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010011110000111101)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010011110000111110) && ({row_reg, col_reg}<18'b010011110001000000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011110001000000)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010011110001000001) && ({row_reg, col_reg}<18'b010011110001000011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010011110001000011) && ({row_reg, col_reg}<18'b010011110001000101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010011110001000101) && ({row_reg, col_reg}<18'b010011110001001000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011110001001000)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==18'b010011110001001001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010011110001001010)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010011110001001011) && ({row_reg, col_reg}<18'b010011110001001101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011110001001101)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==18'b010011110001001110)) color_data = 12'b011001111000;
		if(({row_reg, col_reg}==18'b010011110001001111)) color_data = 12'b010101111000;
		if(({row_reg, col_reg}==18'b010011110001010000)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}>=18'b010011110001010001) && ({row_reg, col_reg}<18'b010011110001010100)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010011110001010100)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b010011110001010101)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b010011110001010110)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}>=18'b010011110001010111) && ({row_reg, col_reg}<18'b010011110001011001)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b010011110001011001)) color_data = 12'b011011001110;
		if(({row_reg, col_reg}==18'b010011110001011010)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010011110001011011) && ({row_reg, col_reg}<18'b010011110001011111)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010011110001011111) && ({row_reg, col_reg}<18'b010011110001100010)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010011110001100010)) color_data = 12'b100011011111;
		if(({row_reg, col_reg}==18'b010011110001100011)) color_data = 12'b001110001011;
		if(({row_reg, col_reg}==18'b010011110001100100)) color_data = 12'b001101111011;
		if(({row_reg, col_reg}>=18'b010011110001100101) && ({row_reg, col_reg}<18'b010011110001101001)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010011110001101001)) color_data = 12'b010010001011;
		if(({row_reg, col_reg}==18'b010011110001101010)) color_data = 12'b010001111010;
		if(({row_reg, col_reg}==18'b010011110001101011)) color_data = 12'b010101111001;
		if(({row_reg, col_reg}==18'b010011110001101100)) color_data = 12'b100010011010;
		if(({row_reg, col_reg}==18'b010011110001101101)) color_data = 12'b101010111100;
		if(({row_reg, col_reg}==18'b010011110001101110)) color_data = 12'b101010101100;
		if(({row_reg, col_reg}>=18'b010011110001101111) && ({row_reg, col_reg}<18'b010011110001110010)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}>=18'b010011110001110010) && ({row_reg, col_reg}<18'b010011110001110100)) color_data = 12'b101010101100;
		if(({row_reg, col_reg}>=18'b010011110001110100) && ({row_reg, col_reg}<18'b010011110001110111)) color_data = 12'b101010101101;
		if(({row_reg, col_reg}==18'b010011110001110111)) color_data = 12'b101010111100;
		if(({row_reg, col_reg}==18'b010011110001111000)) color_data = 12'b101010101100;
		if(({row_reg, col_reg}==18'b010011110001111001)) color_data = 12'b101010111100;
		if(({row_reg, col_reg}==18'b010011110001111010)) color_data = 12'b101010101100;
		if(({row_reg, col_reg}==18'b010011110001111011)) color_data = 12'b101010111100;
		if(({row_reg, col_reg}==18'b010011110001111100)) color_data = 12'b101010101100;
		if(({row_reg, col_reg}==18'b010011110001111101)) color_data = 12'b101010111100;
		if(({row_reg, col_reg}==18'b010011110001111110)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b010011110001111111)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}>=18'b010011110010000000) && ({row_reg, col_reg}<18'b010011110010000011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011110010000011)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010011110010000100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010011110010000101)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b010011110010000110) && ({row_reg, col_reg}<18'b010011110010001100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010011110010001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010011110010001101)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010011110010001110)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010011110010001111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010011110010010000) && ({row_reg, col_reg}<18'b010011110010010010)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010011110010010010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010011110010010011) && ({row_reg, col_reg}<18'b010011110010011011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011110010011011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010011110010011100) && ({row_reg, col_reg}<18'b010011110010101010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010011110010101010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010011110010101011) && ({row_reg, col_reg}<18'b010011110010110011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011110010110011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010011110010110100) && ({row_reg, col_reg}<18'b010011110010111000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010011110010111000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b010011110010111001) && ({row_reg, col_reg}<18'b010011110010111111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011110010111111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010011110011000000) && ({row_reg, col_reg}<18'b010011110011000101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010011110011000101) && ({row_reg, col_reg}<18'b010011110011000111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010011110011000111) && ({row_reg, col_reg}<18'b010011110011001001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010011110011001001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010011110011001010) && ({row_reg, col_reg}<18'b010011110011001100)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010011110011001100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010011110011001101)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b010011110011001110) && ({row_reg, col_reg}<18'b010011110011010000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010011110011010000)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010011110011010001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010011110011010010)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b010011110011010011) && ({row_reg, col_reg}<18'b010011110011011110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010011110011011110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010011110011011111) && ({row_reg, col_reg}<18'b010011110011100011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011110011100011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010011110011100100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010011110011100101) && ({row_reg, col_reg}<18'b010011110011110011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011110011110011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010011110011110100) && ({row_reg, col_reg}<18'b010011110011111000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011110011111000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010011110011111001) && ({row_reg, col_reg}<18'b010011110011111110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011110011111110)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}==18'b010011110011111111)) color_data = 12'b011001101000;
		if(({row_reg, col_reg}>=18'b010011110100000000) && ({row_reg, col_reg}<18'b010011110100000010)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}>=18'b010011110100000010) && ({row_reg, col_reg}<18'b010011110100000100)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}>=18'b010011110100000100) && ({row_reg, col_reg}<18'b010011110100000110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010011110100000110) && ({row_reg, col_reg}<18'b010011110100001000)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b010011110100001000) && ({row_reg, col_reg}<18'b010011110100001010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010011110100001010) && ({row_reg, col_reg}<18'b010011110100001100)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b010011110100001100) && ({row_reg, col_reg}<18'b010011111000000100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010011111000000100) && ({row_reg, col_reg}<18'b010011111000000111)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010011111000000111) && ({row_reg, col_reg}<18'b010011111000001001)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}==18'b010011111000001001)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010011111000001010) && ({row_reg, col_reg}<18'b010011111000001100)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}>=18'b010011111000001100) && ({row_reg, col_reg}<18'b010011111000010000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010011111000010000)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b010011111000010001)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==18'b010011111000010010)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}>=18'b010011111000010011) && ({row_reg, col_reg}<18'b010011111000010101)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b010011111000010101) && ({row_reg, col_reg}<18'b010011111000010111)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010011111000010111)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}==18'b010011111000011000)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b010011111000011001)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b010011111000011010)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b010011111000011011)) color_data = 12'b011011001110;
		if(({row_reg, col_reg}>=18'b010011111000011100) && ({row_reg, col_reg}<18'b010011111000100000)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010011111000100000)) color_data = 12'b010110111101;
		if(({row_reg, col_reg}==18'b010011111000100001)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}>=18'b010011111000100010) && ({row_reg, col_reg}<18'b010011111000100100)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b010011111000100100)) color_data = 12'b010110001011;
		if(({row_reg, col_reg}==18'b010011111000100101)) color_data = 12'b010101111000;
		if(({row_reg, col_reg}==18'b010011111000100110)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}==18'b010011111000100111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010011111000101000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011111000101001)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010011111000101010) && ({row_reg, col_reg}<18'b010011111000101100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010011111000101100) && ({row_reg, col_reg}<18'b010011111000101111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011111000101111)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010011111000110000) && ({row_reg, col_reg}<18'b010011111000110011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011111000110011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010011111000110100) && ({row_reg, col_reg}<18'b010011111000111000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010011111000111000) && ({row_reg, col_reg}<18'b010011111000111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010011111000111100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010011111000111101) && ({row_reg, col_reg}<18'b010011111001000011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011111001000011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010011111001000100)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==18'b010011111001000101)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}>=18'b010011111001000110) && ({row_reg, col_reg}<18'b010011111001001001)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010011111001001001) && ({row_reg, col_reg}<18'b010011111001001011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010011111001001011) && ({row_reg, col_reg}<18'b010011111001001101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011111001001101)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}==18'b010011111001001110)) color_data = 12'b011001111000;
		if(({row_reg, col_reg}==18'b010011111001001111)) color_data = 12'b010101111000;
		if(({row_reg, col_reg}>=18'b010011111001010000) && ({row_reg, col_reg}<18'b010011111001010011)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010011111001010011)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010011111001010100)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b010011111001010101)) color_data = 12'b001110011100;
		if(({row_reg, col_reg}==18'b010011111001010110)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}>=18'b010011111001010111) && ({row_reg, col_reg}<18'b010011111001011001)) color_data = 12'b001010011011;
		if(({row_reg, col_reg}==18'b010011111001011001)) color_data = 12'b011011011111;
		if(({row_reg, col_reg}>=18'b010011111001011010) && ({row_reg, col_reg}<18'b010011111001011100)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010011111001011100)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010011111001011101)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010011111001011110) && ({row_reg, col_reg}<18'b010011111001100001)) color_data = 12'b011111101111;
		if(({row_reg, col_reg}>=18'b010011111001100001) && ({row_reg, col_reg}<18'b010011111001100011)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}==18'b010011111001100011)) color_data = 12'b001110011011;
		if(({row_reg, col_reg}>=18'b010011111001100100) && ({row_reg, col_reg}<18'b010011111001101000)) color_data = 12'b010010001100;
		if(({row_reg, col_reg}==18'b010011111001101000)) color_data = 12'b001101111011;
		if(({row_reg, col_reg}==18'b010011111001101001)) color_data = 12'b010001111011;
		if(({row_reg, col_reg}==18'b010011111001101010)) color_data = 12'b010001111010;
		if(({row_reg, col_reg}==18'b010011111001101011)) color_data = 12'b011010001001;
		if(({row_reg, col_reg}==18'b010011111001101100)) color_data = 12'b100010011011;
		if(({row_reg, col_reg}==18'b010011111001101101)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b010011111001101110)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b010011111001101111)) color_data = 12'b101010101100;
		if(({row_reg, col_reg}>=18'b010011111001110000) && ({row_reg, col_reg}<18'b010011111001110010)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b010011111001110010)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b010011111001110011)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==18'b010011111001110100)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b010011111001110101)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}==18'b010011111001110110)) color_data = 12'b100110101101;
		if(({row_reg, col_reg}>=18'b010011111001110111) && ({row_reg, col_reg}<18'b010011111001111001)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==18'b010011111001111001)) color_data = 12'b100010011100;
		if(({row_reg, col_reg}>=18'b010011111001111010) && ({row_reg, col_reg}<18'b010011111001111100)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}>=18'b010011111001111100) && ({row_reg, col_reg}<18'b010011111001111111)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b010011111001111111)) color_data = 12'b011110001001;
		if(({row_reg, col_reg}==18'b010011111010000000)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010011111010000001) && ({row_reg, col_reg}<18'b010011111010000011)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==18'b010011111010000011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011111010000100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010011111010000101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010011111010000110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010011111010000111) && ({row_reg, col_reg}<18'b010011111010001100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010011111010001100) && ({row_reg, col_reg}<18'b010011111010001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010011111010001110) && ({row_reg, col_reg}<18'b010011111010010000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b010011111010010000) && ({row_reg, col_reg}<18'b010011111010010010)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010011111010010010)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b010011111010010011) && ({row_reg, col_reg}<18'b010011111010011011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011111010011011)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010011111010011100) && ({row_reg, col_reg}<18'b010011111010011110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010011111010011110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010011111010011111) && ({row_reg, col_reg}<18'b010011111010100010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010011111010100010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010011111010100011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010011111010100100) && ({row_reg, col_reg}<18'b010011111010100110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010011111010100110) && ({row_reg, col_reg}<18'b010011111010101001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010011111010101001) && ({row_reg, col_reg}<18'b010011111010101011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010011111010101011) && ({row_reg, col_reg}<18'b010011111010110011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011111010110011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010011111010110100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010011111010110101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010011111010110110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010011111010110111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010011111010111000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b010011111010111001) && ({row_reg, col_reg}<18'b010011111010111011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011111010111011)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010011111010111100) && ({row_reg, col_reg}<18'b010011111011000101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010011111011000101) && ({row_reg, col_reg}<18'b010011111011000111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010011111011000111) && ({row_reg, col_reg}<18'b010011111011001001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010011111011001001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010011111011001010) && ({row_reg, col_reg}<18'b010011111011001110)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010011111011001110)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==18'b010011111011001111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010011111011010000)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b010011111011010001) && ({row_reg, col_reg}<18'b010011111011010011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010011111011010011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010011111011010100) && ({row_reg, col_reg}<18'b010011111011011110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010011111011011110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010011111011011111) && ({row_reg, col_reg}<18'b010011111011110011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010011111011110011) && ({row_reg, col_reg}<18'b010011111011110101)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010011111011110101) && ({row_reg, col_reg}<18'b010011111011110111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010011111011110111) && ({row_reg, col_reg}<18'b010011111011111010)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010011111011111010) && ({row_reg, col_reg}<18'b010011111011111101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010011111011111101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010011111011111110) && ({row_reg, col_reg}<18'b010011111100000000)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}==18'b010011111100000000)) color_data = 12'b100010111100;
		if(({row_reg, col_reg}==18'b010011111100000001)) color_data = 12'b100010111101;
		if(({row_reg, col_reg}==18'b010011111100000010)) color_data = 12'b011110111101;
		if(({row_reg, col_reg}==18'b010011111100000011)) color_data = 12'b011110111110;
		if(({row_reg, col_reg}==18'b010011111100000100)) color_data = 12'b011110111111;
		if(({row_reg, col_reg}==18'b010011111100000101)) color_data = 12'b011010111111;
		if(({row_reg, col_reg}>=18'b010011111100000110) && ({row_reg, col_reg}<18'b010011111100001000)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b010011111100001000) && ({row_reg, col_reg}<18'b010011111100001010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010011111100001010) && ({row_reg, col_reg}<18'b010011111100001100)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b010011111100001100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010011111100001101)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b010011111100001110) && ({row_reg, col_reg}<18'b010100000000000100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010100000000000100)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010100000000000101) && ({row_reg, col_reg}<18'b010100000000000111)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}>=18'b010100000000000111) && ({row_reg, col_reg}<18'b010100000000001011)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010100000000001011) && ({row_reg, col_reg}<18'b010100000000001110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010100000000001110)) color_data = 12'b011110111110;
		if(({row_reg, col_reg}>=18'b010100000000001111) && ({row_reg, col_reg}<18'b010100000000010001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010100000000010001)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b010100000000010010)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}>=18'b010100000000010011) && ({row_reg, col_reg}<18'b010100000000011001)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b010100000000011001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010100000000011010)) color_data = 12'b010110101101;
		if(({row_reg, col_reg}==18'b010100000000011011)) color_data = 12'b100011011111;
		if(({row_reg, col_reg}==18'b010100000000011100)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010100000000011101)) color_data = 12'b100011101110;
		if(({row_reg, col_reg}==18'b010100000000011110)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010100000000011111)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010100000000100000) && ({row_reg, col_reg}<18'b010100000000100010)) color_data = 12'b011111101111;
		if(({row_reg, col_reg}==18'b010100000000100010)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010100000000100011)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b010100000000100100)) color_data = 12'b100111001101;
		if(({row_reg, col_reg}==18'b010100000000100101)) color_data = 12'b011010001000;
		if(({row_reg, col_reg}==18'b010100000000100110)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==18'b010100000000100111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010100000000101000)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==18'b010100000000101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010100000000101010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010100000000101011) && ({row_reg, col_reg}<18'b010100000000101101)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010100000000101101) && ({row_reg, col_reg}<18'b010100000000110011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010100000000110011) && ({row_reg, col_reg}<18'b010100000000110110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010100000000110110)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010100000000110111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010100000000111000) && ({row_reg, col_reg}<18'b010100000000111011)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010100000000111011) && ({row_reg, col_reg}<18'b010100000000111110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010100000000111110) && ({row_reg, col_reg}<18'b010100000001000001)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010100000001000001) && ({row_reg, col_reg}<18'b010100000001000110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010100000001000110) && ({row_reg, col_reg}<18'b010100000001001000)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010100000001001000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010100000001001001) && ({row_reg, col_reg}<18'b010100000001001011)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010100000001001011) && ({row_reg, col_reg}<18'b010100000001001101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100000001001101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010100000001001110)) color_data = 12'b011001111000;
		if(({row_reg, col_reg}==18'b010100000001001111)) color_data = 12'b010101111000;
		if(({row_reg, col_reg}==18'b010100000001010000)) color_data = 12'b001101111011;
		if(({row_reg, col_reg}==18'b010100000001010001)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}>=18'b010100000001010010) && ({row_reg, col_reg}<18'b010100000001010100)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010100000001010100)) color_data = 12'b010110101110;
		if(({row_reg, col_reg}==18'b010100000001010101)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}>=18'b010100000001010110) && ({row_reg, col_reg}<18'b010100000001011000)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010100000001011000)) color_data = 12'b011111101110;
		if(({row_reg, col_reg}>=18'b010100000001011001) && ({row_reg, col_reg}<18'b010100000001011101)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010100000001011101)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010100000001011110)) color_data = 12'b010010101100;
		if(({row_reg, col_reg}==18'b010100000001011111)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b010100000001100000)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b010100000001100001)) color_data = 12'b001110011100;
		if(({row_reg, col_reg}==18'b010100000001100010)) color_data = 12'b001110101100;
		if(({row_reg, col_reg}>=18'b010100000001100011) && ({row_reg, col_reg}<18'b010100000001100101)) color_data = 12'b011111101111;
		if(({row_reg, col_reg}>=18'b010100000001100101) && ({row_reg, col_reg}<18'b010100000001100111)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010100000001100111)) color_data = 12'b100011001101;
		if(({row_reg, col_reg}>=18'b010100000001101000) && ({row_reg, col_reg}<18'b010100000001101010)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}==18'b010100000001101010)) color_data = 12'b100110011011;
		if(({row_reg, col_reg}==18'b010100000001101011)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}==18'b010100000001101100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010100000001101101) && ({row_reg, col_reg}<18'b010100000001110000)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b010100000001110000)) color_data = 12'b100010101010;
		if(({row_reg, col_reg}==18'b010100000001110001)) color_data = 12'b011010011001;
		if(({row_reg, col_reg}==18'b010100000001110010)) color_data = 12'b010101111001;
		if(({row_reg, col_reg}==18'b010100000001110011)) color_data = 12'b010101111011;
		if(({row_reg, col_reg}==18'b010100000001110100)) color_data = 12'b010001111100;
		if(({row_reg, col_reg}>=18'b010100000001110101) && ({row_reg, col_reg}<18'b010100000001110111)) color_data = 12'b010001111101;
		if(({row_reg, col_reg}==18'b010100000001110111)) color_data = 12'b010001111100;
		if(({row_reg, col_reg}==18'b010100000001111000)) color_data = 12'b010001111011;
		if(({row_reg, col_reg}>=18'b010100000001111001) && ({row_reg, col_reg}<18'b010100000001111011)) color_data = 12'b010010001011;
		if(({row_reg, col_reg}==18'b010100000001111011)) color_data = 12'b001101111011;
		if(({row_reg, col_reg}>=18'b010100000001111100) && ({row_reg, col_reg}<18'b010100000001111110)) color_data = 12'b010001111010;
		if(({row_reg, col_reg}==18'b010100000001111110)) color_data = 12'b010110001010;
		if(({row_reg, col_reg}==18'b010100000001111111)) color_data = 12'b010101111010;
		if(({row_reg, col_reg}==18'b010100000010000000)) color_data = 12'b010101110111;
		if(({row_reg, col_reg}>=18'b010100000010000001) && ({row_reg, col_reg}<18'b010100000010000011)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}>=18'b010100000010000011) && ({row_reg, col_reg}<18'b010100000010000101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100000010000101)) color_data = 12'b100001110101;
		if(({row_reg, col_reg}==18'b010100000010000110)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}>=18'b010100000010000111) && ({row_reg, col_reg}<18'b010100000010001001)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010100000010001001) && ({row_reg, col_reg}<18'b010100000010001011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010100000010001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010100000010001100) && ({row_reg, col_reg}<18'b010100000010001110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010100000010001110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010100000010001111)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}==18'b010100000010010000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010100000010010001)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010100000010010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010100000010010011) && ({row_reg, col_reg}<18'b010100000010100000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010100000010100000) && ({row_reg, col_reg}<18'b010100000010100010)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010100000010100010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010100000010100011) && ({row_reg, col_reg}<18'b010100000010100101)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==18'b010100000010100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010100000010100110) && ({row_reg, col_reg}<18'b010100000010101000)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010100000010101000) && ({row_reg, col_reg}<18'b010100000010101011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100000010101011)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010100000010101100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010100000010101101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100000010101110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010100000010101111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100000010110000)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}>=18'b010100000010110001) && ({row_reg, col_reg}<18'b010100000010110011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100000010110011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010100000010110100)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==18'b010100000010110101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010100000010110110)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010100000010110111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010100000010111000)) color_data = 12'b100110001001;
		if(({row_reg, col_reg}>=18'b010100000010111001) && ({row_reg, col_reg}<18'b010100000011000111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100000011000111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010100000011001000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010100000011001001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010100000011001010)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010100000011001011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010100000011001100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010100000011001101)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010100000011001110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010100000011001111)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010100000011010000) && ({row_reg, col_reg}<18'b010100000011011111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010100000011011111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010100000011100000) && ({row_reg, col_reg}<18'b010100000011110000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010100000011110000) && ({row_reg, col_reg}<18'b010100000011110010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010100000011110010) && ({row_reg, col_reg}<18'b010100000011111000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100000011111000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010100000011111001) && ({row_reg, col_reg}<18'b010100000011111100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100000011111100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010100000011111101)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}==18'b010100000011111110)) color_data = 12'b010101110110;
		if(({row_reg, col_reg}==18'b010100000011111111)) color_data = 12'b010101110111;
		if(({row_reg, col_reg}==18'b010100000100000000)) color_data = 12'b100011011100;
		if(({row_reg, col_reg}==18'b010100000100000001)) color_data = 12'b100111101110;
		if(({row_reg, col_reg}>=18'b010100000100000010) && ({row_reg, col_reg}<18'b010100000100000100)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b010100000100000100)) color_data = 12'b100011011111;
		if(({row_reg, col_reg}==18'b010100000100000101)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}>=18'b010100000100000110) && ({row_reg, col_reg}<18'b010100000100001001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010100000100001001) && ({row_reg, col_reg}<18'b010100000100001100)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b010100000100001100) && ({row_reg, col_reg}<18'b010100001000001011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010100001000001011) && ({row_reg, col_reg}<18'b010100001000001101)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}>=18'b010100001000001101) && ({row_reg, col_reg}<18'b010100001000010001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010100001000010001)) color_data = 12'b011110111111;
		if(({row_reg, col_reg}==18'b010100001000010010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010100001000010011) && ({row_reg, col_reg}<18'b010100001000011001)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b010100001000011001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010100001000011010)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}==18'b010100001000011011)) color_data = 12'b011111011110;
		if(({row_reg, col_reg}==18'b010100001000011100)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010100001000011101) && ({row_reg, col_reg}<18'b010100001000100011)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010100001000100011)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}==18'b010100001000100100)) color_data = 12'b100111011101;
		if(({row_reg, col_reg}==18'b010100001000100101)) color_data = 12'b010101111000;
		if(({row_reg, col_reg}==18'b010100001000100110)) color_data = 12'b010101100110;
		if(({row_reg, col_reg}>=18'b010100001000100111) && ({row_reg, col_reg}<18'b010100001000101001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010100001000101001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010100001000101010) && ({row_reg, col_reg}<18'b010100001000101101)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010100001000101101) && ({row_reg, col_reg}<18'b010100001000101111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100001000101111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010100001000110000) && ({row_reg, col_reg}<18'b010100001000110010)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010100001000110010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010100001000110011) && ({row_reg, col_reg}<18'b010100001000110110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010100001000110110)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b010100001000110111) && ({row_reg, col_reg}<18'b010100001000111010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010100001000111010) && ({row_reg, col_reg}<18'b010100001001000000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100001001000000)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}>=18'b010100001001000001) && ({row_reg, col_reg}<18'b010100001001000111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100001001000111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010100001001001000) && ({row_reg, col_reg}<18'b010100001001001010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100001001001010)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010100001001001011) && ({row_reg, col_reg}<18'b010100001001001101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100001001001101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010100001001001110)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==18'b010100001001001111)) color_data = 12'b010101111000;
		if(({row_reg, col_reg}==18'b010100001001010000)) color_data = 12'b001110001011;
		if(({row_reg, col_reg}==18'b010100001001010001)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010100001001010010)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010100001001010011)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010100001001010100)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==18'b010100001001010101)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010100001001010110) && ({row_reg, col_reg}<18'b010100001001011010)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010100001001011010)) color_data = 12'b011111111110;
		if(({row_reg, col_reg}==18'b010100001001011011)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010100001001011100)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010100001001011101)) color_data = 12'b011111101111;
		if(({row_reg, col_reg}==18'b010100001001011110)) color_data = 12'b001110011100;
		if(({row_reg, col_reg}==18'b010100001001011111)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b010100001001100000)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b010100001001100001)) color_data = 12'b000110001011;
		if(({row_reg, col_reg}==18'b010100001001100010)) color_data = 12'b001110011100;
		if(({row_reg, col_reg}>=18'b010100001001100011) && ({row_reg, col_reg}<18'b010100001001100101)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010100001001100101)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010100001001100110)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b010100001001100111)) color_data = 12'b100111001101;
		if(({row_reg, col_reg}==18'b010100001001101000)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}==18'b010100001001101001)) color_data = 12'b100010011010;
		if(({row_reg, col_reg}==18'b010100001001101010)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}==18'b010100001001101011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010100001001101100)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}>=18'b010100001001101101) && ({row_reg, col_reg}<18'b010100001001101111)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b010100001001101111)) color_data = 12'b101010111100;
		if(({row_reg, col_reg}==18'b010100001001110000)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b010100001001110001)) color_data = 12'b011010001001;
		if(({row_reg, col_reg}==18'b010100001001110010)) color_data = 12'b010001101001;
		if(({row_reg, col_reg}==18'b010100001001110011)) color_data = 12'b010001111011;
		if(({row_reg, col_reg}==18'b010100001001110100)) color_data = 12'b010001111100;
		if(({row_reg, col_reg}==18'b010100001001110101)) color_data = 12'b010001111101;
		if(({row_reg, col_reg}>=18'b010100001001110110) && ({row_reg, col_reg}<18'b010100001001111000)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010100001001111000)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}>=18'b010100001001111001) && ({row_reg, col_reg}<18'b010100001001111101)) color_data = 12'b001101111011;
		if(({row_reg, col_reg}==18'b010100001001111101)) color_data = 12'b010001111011;
		if(({row_reg, col_reg}==18'b010100001001111110)) color_data = 12'b010001111010;
		if(({row_reg, col_reg}==18'b010100001001111111)) color_data = 12'b010001111001;
		if(({row_reg, col_reg}==18'b010100001010000000)) color_data = 12'b010101100111;
		if(({row_reg, col_reg}==18'b010100001010000001)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==18'b010100001010000010)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}==18'b010100001010000011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010100001010000100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100001010000101)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010100001010000110)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==18'b010100001010000111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010100001010001000) && ({row_reg, col_reg}<18'b010100001010001010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010100001010001010) && ({row_reg, col_reg}<18'b010100001010010001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010100001010010001)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010100001010010010)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010100001010010011) && ({row_reg, col_reg}<18'b010100001010100000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100001010100000)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010100001010100001) && ({row_reg, col_reg}<18'b010100001010110011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100001010110011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010100001010110100) && ({row_reg, col_reg}<18'b010100001010110110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010100001010110110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010100001010110111)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==18'b010100001010111000)) color_data = 12'b100110001001;
		if(({row_reg, col_reg}==18'b010100001010111001)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010100001010111010) && ({row_reg, col_reg}<18'b010100001011000001)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100001011000001)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010100001011000010) && ({row_reg, col_reg}<18'b010100001011000111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100001011000111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010100001011001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010100001011001001) && ({row_reg, col_reg}<18'b010100001011011110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010100001011011110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010100001011011111) && ({row_reg, col_reg}<18'b010100001011110000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100001011110000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010100001011110001) && ({row_reg, col_reg}<18'b010100001011111101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100001011111101)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}==18'b010100001011111110)) color_data = 12'b010101110110;
		if(({row_reg, col_reg}==18'b010100001011111111)) color_data = 12'b011010000111;
		if(({row_reg, col_reg}==18'b010100001100000000)) color_data = 12'b100111101110;
		if(({row_reg, col_reg}>=18'b010100001100000001) && ({row_reg, col_reg}<18'b010100001100000100)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}==18'b010100001100000100)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b010100001100000101)) color_data = 12'b011110111110;
		if(({row_reg, col_reg}>=18'b010100001100000110) && ({row_reg, col_reg}<18'b010100001100001000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010100001100001000)) color_data = 12'b011110111110;

		if(({row_reg, col_reg}>=18'b010100001100001001) && ({row_reg, col_reg}<18'b010100010000000110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010100010000000110) && ({row_reg, col_reg}<18'b010100010000001001)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010100010000001001) && ({row_reg, col_reg}<18'b010100010000001110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010100010000001110)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}>=18'b010100010000001111) && ({row_reg, col_reg}<18'b010100010000010001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010100010000010001)) color_data = 12'b011110111110;
		if(({row_reg, col_reg}>=18'b010100010000010010) && ({row_reg, col_reg}<18'b010100010000010101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010100010000010101) && ({row_reg, col_reg}<18'b010100010000010111)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b010100010000010111) && ({row_reg, col_reg}<18'b010100010000011001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010100010000011001)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==18'b010100010000011010)) color_data = 12'b010110111101;
		if(({row_reg, col_reg}==18'b010100010000011011)) color_data = 12'b011111011110;
		if(({row_reg, col_reg}>=18'b010100010000011100) && ({row_reg, col_reg}<18'b010100010000011110)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010100010000011110) && ({row_reg, col_reg}<18'b010100010000100011)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010100010000100011)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010100010000100100)) color_data = 12'b100111011110;
		if(({row_reg, col_reg}==18'b010100010000100101)) color_data = 12'b010110001001;
		if(({row_reg, col_reg}==18'b010100010000100110)) color_data = 12'b010101110111;
		if(({row_reg, col_reg}==18'b010100010000100111)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==18'b010100010000101000)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}==18'b010100010000101001)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==18'b010100010000101010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010100010000101011) && ({row_reg, col_reg}<18'b010100010000101101)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010100010000101101) && ({row_reg, col_reg}<18'b010100010000101111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100010000101111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010100010000110000) && ({row_reg, col_reg}<18'b010100010000110010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010100010000110010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100010000110011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010100010000110100) && ({row_reg, col_reg}<18'b010100010000110111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010100010000110111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010100010000111000) && ({row_reg, col_reg}<18'b010100010001001011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100010001001011)) color_data = 12'b100001100110;
		if(({row_reg, col_reg}==18'b010100010001001100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100010001001101)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010100010001001110)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==18'b010100010001001111)) color_data = 12'b010101111000;
		if(({row_reg, col_reg}==18'b010100010001010000)) color_data = 12'b001101111011;
		if(({row_reg, col_reg}>=18'b010100010001010001) && ({row_reg, col_reg}<18'b010100010001010011)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010100010001010011)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010100010001010100)) color_data = 12'b010110101101;
		if(({row_reg, col_reg}==18'b010100010001010101)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010100010001010110) && ({row_reg, col_reg}<18'b010100010001011100)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010100010001011100)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010100010001011101)) color_data = 12'b011111101111;
		if(({row_reg, col_reg}==18'b010100010001011110)) color_data = 12'b010010101100;
		if(({row_reg, col_reg}==18'b010100010001011111)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b010100010001100000)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b010100010001100001)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b010100010001100010)) color_data = 12'b001110011100;
		if(({row_reg, col_reg}>=18'b010100010001100011) && ({row_reg, col_reg}<18'b010100010001100101)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010100010001100101)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}==18'b010100010001100110)) color_data = 12'b101011101111;
		if(({row_reg, col_reg}==18'b010100010001100111)) color_data = 12'b101011001100;
		if(({row_reg, col_reg}==18'b010100010001101000)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}>=18'b010100010001101001) && ({row_reg, col_reg}<18'b010100010001101011)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010100010001101011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010100010001101100)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==18'b010100010001101101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010100010001101110)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b010100010001101111)) color_data = 12'b101010111100;
		if(({row_reg, col_reg}==18'b010100010001110000)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==18'b010100010001110001)) color_data = 12'b011110001011;
		if(({row_reg, col_reg}==18'b010100010001110010)) color_data = 12'b010101111010;
		if(({row_reg, col_reg}==18'b010100010001110011)) color_data = 12'b010101111011;
		if(({row_reg, col_reg}==18'b010100010001110100)) color_data = 12'b010001111100;
		if(({row_reg, col_reg}==18'b010100010001110101)) color_data = 12'b010001111101;
		if(({row_reg, col_reg}>=18'b010100010001110110) && ({row_reg, col_reg}<18'b010100010001111011)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010100010001111011)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b010100010001111100) && ({row_reg, col_reg}<18'b010100010001111110)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010100010001111110)) color_data = 12'b010001111011;
		if(({row_reg, col_reg}==18'b010100010001111111)) color_data = 12'b010001111010;
		if(({row_reg, col_reg}>=18'b010100010010000000) && ({row_reg, col_reg}<18'b010100010010000010)) color_data = 12'b010101111000;
		if(({row_reg, col_reg}>=18'b010100010010000010) && ({row_reg, col_reg}<18'b010100010010000100)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}>=18'b010100010010000100) && ({row_reg, col_reg}<18'b010100010010001000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100010010001000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010100010010001001) && ({row_reg, col_reg}<18'b010100010010001100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010100010010001100)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b010100010010001101) && ({row_reg, col_reg}<18'b010100010010010010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010100010010010010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010100010010010011) && ({row_reg, col_reg}<18'b010100010010110000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010100010010110000) && ({row_reg, col_reg}<18'b010100010010110011)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==18'b010100010010110011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010100010010110100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010100010010110101) && ({row_reg, col_reg}<18'b010100010010110111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010100010010110111)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==18'b010100010010111000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b010100010010111001) && ({row_reg, col_reg}<18'b010100010010111011)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010100010010111011) && ({row_reg, col_reg}<18'b010100010010111101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100010010111101)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010100010010111110) && ({row_reg, col_reg}<18'b010100010011000101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100010011000101)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010100010011000110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010100010011000111) && ({row_reg, col_reg}<18'b010100010011011110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010100010011011110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010100010011011111) && ({row_reg, col_reg}<18'b010100010011111000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100010011111000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010100010011111001) && ({row_reg, col_reg}<18'b010100010011111101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100010011111101)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010100010011111110)) color_data = 12'b010101100110;
		if(({row_reg, col_reg}==18'b010100010011111111)) color_data = 12'b011010000111;
		if(({row_reg, col_reg}==18'b010100010100000000)) color_data = 12'b100111011110;
		if(({row_reg, col_reg}==18'b010100010100000001)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}>=18'b010100010100000010) && ({row_reg, col_reg}<18'b010100010100000100)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010100010100000100)) color_data = 12'b100011011111;
		if(({row_reg, col_reg}==18'b010100010100000101)) color_data = 12'b011110111110;
		if(({row_reg, col_reg}>=18'b010100010100000110) && ({row_reg, col_reg}<18'b010100010100001010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010100010100001010) && ({row_reg, col_reg}<18'b010100010100001101)) color_data = 12'b011010101101;

		if(({row_reg, col_reg}>=18'b010100010100001101) && ({row_reg, col_reg}<18'b010100011000000001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010100011000000001)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010100011000000010) && ({row_reg, col_reg}<18'b010100011000000110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010100011000000110) && ({row_reg, col_reg}<18'b010100011000001000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010100011000001000) && ({row_reg, col_reg}<18'b010100011000001010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010100011000001010)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}>=18'b010100011000001011) && ({row_reg, col_reg}<18'b010100011000010110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010100011000010110)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==18'b010100011000010111)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}==18'b010100011000011000)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}==18'b010100011000011001)) color_data = 12'b010110111101;
		if(({row_reg, col_reg}==18'b010100011000011010)) color_data = 12'b010110111100;
		if(({row_reg, col_reg}==18'b010100011000011011)) color_data = 12'b011111101110;
		if(({row_reg, col_reg}==18'b010100011000011100)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010100011000011101) && ({row_reg, col_reg}<18'b010100011000100011)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010100011000100011)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010100011000100100)) color_data = 12'b100011011101;
		if(({row_reg, col_reg}==18'b010100011000100101)) color_data = 12'b010110001001;
		if(({row_reg, col_reg}==18'b010100011000100110)) color_data = 12'b001101100110;
		if(({row_reg, col_reg}==18'b010100011000100111)) color_data = 12'b010001100111;
		if(({row_reg, col_reg}==18'b010100011000101000)) color_data = 12'b010101110111;
		if(({row_reg, col_reg}>=18'b010100011000101001) && ({row_reg, col_reg}<18'b010100011000101011)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}==18'b010100011000101011)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010100011000101100) && ({row_reg, col_reg}<18'b010100011000101111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100011000101111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010100011000110000) && ({row_reg, col_reg}<18'b010100011000110010)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}==18'b010100011000110010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010100011000110011) && ({row_reg, col_reg}<18'b010100011000111000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010100011000111000) && ({row_reg, col_reg}<18'b010100011000111010)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010100011000111010) && ({row_reg, col_reg}<18'b010100011000111111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100011000111111)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010100011001000000) && ({row_reg, col_reg}<18'b010100011001000010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010100011001000010) && ({row_reg, col_reg}<18'b010100011001000100)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010100011001000100) && ({row_reg, col_reg}<18'b010100011001001110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100011001001110)) color_data = 12'b010101110111;
		if(({row_reg, col_reg}==18'b010100011001001111)) color_data = 12'b010101111000;
		if(({row_reg, col_reg}==18'b010100011001010000)) color_data = 12'b010010001100;
		if(({row_reg, col_reg}==18'b010100011001010001)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010100011001010010)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010100011001010011)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010100011001010100)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}>=18'b010100011001010101) && ({row_reg, col_reg}<18'b010100011001011011)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010100011001011011)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010100011001011100)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010100011001011101)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010100011001011110)) color_data = 12'b001110011100;
		if(({row_reg, col_reg}==18'b010100011001011111)) color_data = 12'b000101111001;
		if(({row_reg, col_reg}==18'b010100011001100000)) color_data = 12'b001110001011;
		if(({row_reg, col_reg}==18'b010100011001100001)) color_data = 12'b001001111010;
		if(({row_reg, col_reg}==18'b010100011001100010)) color_data = 12'b010010011011;
		if(({row_reg, col_reg}==18'b010100011001100011)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b010100011001100100)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}==18'b010100011001100101)) color_data = 12'b101011101111;
		if(({row_reg, col_reg}==18'b010100011001100110)) color_data = 12'b101111101110;
		if(({row_reg, col_reg}==18'b010100011001100111)) color_data = 12'b101011001100;
		if(({row_reg, col_reg}==18'b010100011001101000)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}>=18'b010100011001101001) && ({row_reg, col_reg}<18'b010100011001101011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010100011001101011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010100011001101100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b010100011001101101) && ({row_reg, col_reg}<18'b010100011001101111)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==18'b010100011001101111)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b010100011001110000)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==18'b010100011001110001)) color_data = 12'b011110001010;
		if(({row_reg, col_reg}==18'b010100011001110010)) color_data = 12'b010101101001;
		if(({row_reg, col_reg}==18'b010100011001110011)) color_data = 12'b010001101010;
		if(({row_reg, col_reg}==18'b010100011001110100)) color_data = 12'b010001111100;
		if(({row_reg, col_reg}>=18'b010100011001110101) && ({row_reg, col_reg}<18'b010100011001110111)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010100011001110111)) color_data = 12'b001001101101;
		if(({row_reg, col_reg}>=18'b010100011001111000) && ({row_reg, col_reg}<18'b010100011001111010)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010100011001111010)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b010100011001111011)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010100011001111100)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b010100011001111101) && ({row_reg, col_reg}<18'b010100011001111111)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010100011001111111)) color_data = 12'b010001111011;
		if(({row_reg, col_reg}>=18'b010100011010000000) && ({row_reg, col_reg}<18'b010100011010000010)) color_data = 12'b010101111001;
		if(({row_reg, col_reg}>=18'b010100011010000010) && ({row_reg, col_reg}<18'b010100011010000100)) color_data = 12'b011001111000;
		if(({row_reg, col_reg}==18'b010100011010000100)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010100011010000101) && ({row_reg, col_reg}<18'b010100011010001001)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010100011010001001) && ({row_reg, col_reg}<18'b010100011010001111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010100011010001111)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}>=18'b010100011010010000) && ({row_reg, col_reg}<18'b010100011010010011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010100011010010011) && ({row_reg, col_reg}<18'b010100011010101101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100011010101101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010100011010101110)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==18'b010100011010101111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100011010110000)) color_data = 12'b100001101000;
		if(({row_reg, col_reg}>=18'b010100011010110001) && ({row_reg, col_reg}<18'b010100011010110011)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==18'b010100011010110011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010100011010110100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010100011010110101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010100011010110110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010100011010110111)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==18'b010100011010111000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010100011010111001)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==18'b010100011010111010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010100011010111011) && ({row_reg, col_reg}<18'b010100011010111110)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010100011010111110) && ({row_reg, col_reg}<18'b010100011011000101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100011011000101)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010100011011000110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010100011011000111) && ({row_reg, col_reg}<18'b010100011011011111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010100011011011111) && ({row_reg, col_reg}<18'b010100011011111101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100011011111101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010100011011111110)) color_data = 12'b010101100110;
		if(({row_reg, col_reg}==18'b010100011011111111)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==18'b010100011100000000)) color_data = 12'b101011101110;
		if(({row_reg, col_reg}==18'b010100011100000001)) color_data = 12'b101011101111;
		if(({row_reg, col_reg}==18'b010100011100000010)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}==18'b010100011100000011)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010100011100000100)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010100011100000101)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}==18'b010100011100000110)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}==18'b010100011100000111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010100011100001000)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}>=18'b010100011100001001) && ({row_reg, col_reg}<18'b010100011100001011)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}>=18'b010100011100001011) && ({row_reg, col_reg}<18'b010100011100001111)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}==18'b010100011100001111)) color_data = 12'b011010101110;

		if(({row_reg, col_reg}>=18'b010100011100010000) && ({row_reg, col_reg}<18'b010100100000000010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010100100000000010) && ({row_reg, col_reg}<18'b010100100000001001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010100100000001001) && ({row_reg, col_reg}<18'b010100100000001011)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}>=18'b010100100000001011) && ({row_reg, col_reg}<18'b010100100000010011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010100100000010011)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010100100000010100) && ({row_reg, col_reg}<18'b010100100000010110)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}==18'b010100100000010110)) color_data = 12'b011110111110;
		if(({row_reg, col_reg}>=18'b010100100000010111) && ({row_reg, col_reg}<18'b010100100000011001)) color_data = 12'b011111001110;
		if(({row_reg, col_reg}==18'b010100100000011001)) color_data = 12'b011111011110;
		if(({row_reg, col_reg}==18'b010100100000011010)) color_data = 12'b011011011101;
		if(({row_reg, col_reg}==18'b010100100000011011)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010100100000011100)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010100100000011101) && ({row_reg, col_reg}<18'b010100100000100000)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010100100000100000)) color_data = 12'b011111111111;
		if(({row_reg, col_reg}>=18'b010100100000100001) && ({row_reg, col_reg}<18'b010100100000100011)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010100100000100011)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010100100000100100)) color_data = 12'b100011011101;
		if(({row_reg, col_reg}==18'b010100100000100101)) color_data = 12'b011111001011;
		if(({row_reg, col_reg}==18'b010100100000100110)) color_data = 12'b011110101010;
		if(({row_reg, col_reg}>=18'b010100100000100111) && ({row_reg, col_reg}<18'b010100100000101001)) color_data = 12'b100010101010;
		if(({row_reg, col_reg}==18'b010100100000101001)) color_data = 12'b011110001001;
		if(({row_reg, col_reg}==18'b010100100000101010)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}>=18'b010100100000101011) && ({row_reg, col_reg}<18'b010100100000101110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010100100000101110) && ({row_reg, col_reg}<18'b010100100000110000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010100100000110000) && ({row_reg, col_reg}<18'b010100100000110010)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}==18'b010100100000110010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010100100000110011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010100100000110100)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010100100000110101) && ({row_reg, col_reg}<18'b010100100000110111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010100100000110111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010100100000111000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010100100000111001) && ({row_reg, col_reg}<18'b010100100000111011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010100100000111011) && ({row_reg, col_reg}<18'b010100100000111111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100100000111111)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010100100001000000) && ({row_reg, col_reg}<18'b010100100001000010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100100001000010)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}==18'b010100100001000011)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010100100001000100) && ({row_reg, col_reg}<18'b010100100001001101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100100001001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010100100001001110)) color_data = 12'b010101110111;
		if(({row_reg, col_reg}==18'b010100100001001111)) color_data = 12'b010101111000;
		if(({row_reg, col_reg}>=18'b010100100001010000) && ({row_reg, col_reg}<18'b010100100001010010)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}>=18'b010100100001010010) && ({row_reg, col_reg}<18'b010100100001010100)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010100100001010100)) color_data = 12'b010010011101;
		if(({row_reg, col_reg}==18'b010100100001010101)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}>=18'b010100100001010110) && ({row_reg, col_reg}<18'b010100100001011011)) color_data = 12'b010110111110;
		if(({row_reg, col_reg}==18'b010100100001011011)) color_data = 12'b011011001110;
		if(({row_reg, col_reg}==18'b010100100001011100)) color_data = 12'b010110111110;
		if(({row_reg, col_reg}==18'b010100100001011101)) color_data = 12'b011011001110;
		if(({row_reg, col_reg}==18'b010100100001011110)) color_data = 12'b010111001101;
		if(({row_reg, col_reg}==18'b010100100001011111)) color_data = 12'b010110111100;
		if(({row_reg, col_reg}>=18'b010100100001100000) && ({row_reg, col_reg}<18'b010100100001100010)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}==18'b010100100001100010)) color_data = 12'b011111001101;
		if(({row_reg, col_reg}==18'b010100100001100011)) color_data = 12'b100011011110;
		if(({row_reg, col_reg}>=18'b010100100001100100) && ({row_reg, col_reg}<18'b010100100001100110)) color_data = 12'b100111001101;
		if(({row_reg, col_reg}==18'b010100100001100110)) color_data = 12'b101011001101;
		if(({row_reg, col_reg}==18'b010100100001100111)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b010100100001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010100100001101001) && ({row_reg, col_reg}<18'b010100100001101100)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010100100001101100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010100100001101101)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b010100100001101110) && ({row_reg, col_reg}<18'b010100100001110000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010100100001110000)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b010100100001110001)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}==18'b010100100001110010)) color_data = 12'b011110001010;
		if(({row_reg, col_reg}==18'b010100100001110011)) color_data = 12'b011110001011;
		if(({row_reg, col_reg}==18'b010100100001110100)) color_data = 12'b011110011101;
		if(({row_reg, col_reg}==18'b010100100001110101)) color_data = 12'b010110011101;
		if(({row_reg, col_reg}==18'b010100100001110110)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010100100001110111)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010100100001111000)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010100100001111001)) color_data = 12'b001010001110;
		if(({row_reg, col_reg}==18'b010100100001111010)) color_data = 12'b001001111111;
		if(({row_reg, col_reg}>=18'b010100100001111011) && ({row_reg, col_reg}<18'b010100100001111101)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b010100100001111101)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010100100001111110)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010100100001111111)) color_data = 12'b001101111011;
		if(({row_reg, col_reg}==18'b010100100010000000)) color_data = 12'b010001111010;
		if(({row_reg, col_reg}==18'b010100100010000001)) color_data = 12'b010101101010;
		if(({row_reg, col_reg}==18'b010100100010000010)) color_data = 12'b010101101001;
		if(({row_reg, col_reg}==18'b010100100010000011)) color_data = 12'b011001101000;
		if(({row_reg, col_reg}==18'b010100100010000100)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}==18'b010100100010000101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010100100010000110) && ({row_reg, col_reg}<18'b010100100010001001)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010100100010001001) && ({row_reg, col_reg}<18'b010100100010001101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010100100010001101)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010100100010001110) && ({row_reg, col_reg}<18'b010100100010010011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010100100010010011) && ({row_reg, col_reg}<18'b010100100010101010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010100100010101010) && ({row_reg, col_reg}<18'b010100100010101101)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010100100010101101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100100010101110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010100100010101111)) color_data = 12'b100101110111;
		if(({row_reg, col_reg}==18'b010100100010110000)) color_data = 12'b100110001001;
		if(({row_reg, col_reg}==18'b010100100010110001)) color_data = 12'b100101111001;
		if(({row_reg, col_reg}>=18'b010100100010110010) && ({row_reg, col_reg}<18'b010100100010110100)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b010100100010110100) && ({row_reg, col_reg}<18'b010100100010110110)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010100100010110110)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==18'b010100100010110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010100100010111000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010100100010111001) && ({row_reg, col_reg}<18'b010100100011000111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100100011000111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010100100011001000) && ({row_reg, col_reg}<18'b010100100011001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010100100011001011) && ({row_reg, col_reg}<18'b010100100011011110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010100100011011110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010100100011011111) && ({row_reg, col_reg}<18'b010100100011110010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010100100011110010) && ({row_reg, col_reg}<18'b010100100011110100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010100100011110100) && ({row_reg, col_reg}<18'b010100100011111101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100100011111101)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010100100011111110)) color_data = 12'b010101110110;
		if(({row_reg, col_reg}==18'b010100100011111111)) color_data = 12'b010101110111;
		if(({row_reg, col_reg}==18'b010100100100000000)) color_data = 12'b100111011110;
		if(({row_reg, col_reg}==18'b010100100100000001)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}>=18'b010100100100000010) && ({row_reg, col_reg}<18'b010100100100000100)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010100100100000100)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010100100100000101)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}==18'b010100100100000110)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}==18'b010100100100000111)) color_data = 12'b011110111110;
		if(({row_reg, col_reg}==18'b010100100100001000)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==18'b010100100100001001)) color_data = 12'b011011001110;
		if(({row_reg, col_reg}==18'b010100100100001010)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}==18'b010100100100001011)) color_data = 12'b011111011110;
		if(({row_reg, col_reg}==18'b010100100100001100)) color_data = 12'b100011011110;
		if(({row_reg, col_reg}==18'b010100100100001101)) color_data = 12'b100011001110;
		if(({row_reg, col_reg}==18'b010100100100001110)) color_data = 12'b011110111110;
		if(({row_reg, col_reg}==18'b010100100100001111)) color_data = 12'b011010111101;

		if(({row_reg, col_reg}>=18'b010100100100010000) && ({row_reg, col_reg}<18'b010100101000000000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010100101000000000) && ({row_reg, col_reg}<18'b010100101000000010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010100101000000010) && ({row_reg, col_reg}<18'b010100101000000110)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}>=18'b010100101000000110) && ({row_reg, col_reg}<18'b010100101000001000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010100101000001000) && ({row_reg, col_reg}<18'b010100101000001011)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010100101000001011) && ({row_reg, col_reg}<18'b010100101000001111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010100101000001111)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b010100101000010000) && ({row_reg, col_reg}<18'b010100101000010100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010100101000010100) && ({row_reg, col_reg}<18'b010100101000010110)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}==18'b010100101000010110)) color_data = 12'b011111001110;
		if(({row_reg, col_reg}==18'b010100101000010111)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}>=18'b010100101000011000) && ({row_reg, col_reg}<18'b010100101000011011)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010100101000011011) && ({row_reg, col_reg}<18'b010100101000100011)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010100101000100011) && ({row_reg, col_reg}<18'b010100101000100101)) color_data = 12'b100011111110;
		if(({row_reg, col_reg}==18'b010100101000100101)) color_data = 12'b100111111110;
		if(({row_reg, col_reg}>=18'b010100101000100110) && ({row_reg, col_reg}<18'b010100101000101000)) color_data = 12'b101111111111;
		if(({row_reg, col_reg}==18'b010100101000101000)) color_data = 12'b110011101110;
		if(({row_reg, col_reg}==18'b010100101000101001)) color_data = 12'b101010111011;
		if(({row_reg, col_reg}==18'b010100101000101010)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==18'b010100101000101011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010100101000101100) && ({row_reg, col_reg}<18'b010100101000101110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100101000101110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010100101000101111)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}==18'b010100101000110000)) color_data = 12'b011001110101;
		if(({row_reg, col_reg}==18'b010100101000110001)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}==18'b010100101000110010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010100101000110011) && ({row_reg, col_reg}<18'b010100101000110101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100101000110101)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010100101000110110) && ({row_reg, col_reg}<18'b010100101000111010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100101000111010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010100101000111011) && ({row_reg, col_reg}<18'b010100101001000001)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010100101001000001) && ({row_reg, col_reg}<18'b010100101001000011)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}==18'b010100101001000011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010100101001000100) && ({row_reg, col_reg}<18'b010100101001001000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100101001001000)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010100101001001001) && ({row_reg, col_reg}<18'b010100101001001101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010100101001001101) && ({row_reg, col_reg}<18'b010100101001001111)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==18'b010100101001001111)) color_data = 12'b010101111000;
		if(({row_reg, col_reg}==18'b010100101001010000)) color_data = 12'b010001111100;
		if(({row_reg, col_reg}==18'b010100101001010001)) color_data = 12'b010001111101;
		if(({row_reg, col_reg}==18'b010100101001010010)) color_data = 12'b010001111110;
		if(({row_reg, col_reg}==18'b010100101001010011)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010100101001010100)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010100101001010101)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010100101001010110)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}>=18'b010100101001010111) && ({row_reg, col_reg}<18'b010100101001011001)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b010100101001011001) && ({row_reg, col_reg}<18'b010100101001011011)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b010100101001011011)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b010100101001011100)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b010100101001011101)) color_data = 12'b001110011100;
		if(({row_reg, col_reg}==18'b010100101001011110)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010100101001011111)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010100101001100000) && ({row_reg, col_reg}<18'b010100101001100010)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}==18'b010100101001100010)) color_data = 12'b101011101111;
		if(({row_reg, col_reg}==18'b010100101001100011)) color_data = 12'b100011001100;
		if(({row_reg, col_reg}==18'b010100101001100100)) color_data = 12'b100010111011;
		if(({row_reg, col_reg}==18'b010100101001100101)) color_data = 12'b100110111011;
		if(({row_reg, col_reg}==18'b010100101001100110)) color_data = 12'b101010111100;
		if(({row_reg, col_reg}==18'b010100101001100111)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}==18'b010100101001101000)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==18'b010100101001101001)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}>=18'b010100101001101010) && ({row_reg, col_reg}<18'b010100101001101100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010100101001101100)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}>=18'b010100101001101101) && ({row_reg, col_reg}<18'b010100101001110000)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010100101001110000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010100101001110001)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==18'b010100101001110010)) color_data = 12'b101010111011;
		if(({row_reg, col_reg}==18'b010100101001110011)) color_data = 12'b100110111100;
		if(({row_reg, col_reg}==18'b010100101001110100)) color_data = 12'b100110111101;
		if(({row_reg, col_reg}==18'b010100101001110101)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b010100101001110110)) color_data = 12'b010010001100;
		if(({row_reg, col_reg}==18'b010100101001110111)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010100101001111000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010100101001111001) && ({row_reg, col_reg}<18'b010100101001111011)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}>=18'b010100101001111011) && ({row_reg, col_reg}<18'b010100101001111101)) color_data = 12'b001001111111;
		if(({row_reg, col_reg}==18'b010100101001111101)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010100101001111110)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010100101001111111)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010100101010000000)) color_data = 12'b010001111100;
		if(({row_reg, col_reg}==18'b010100101010000001)) color_data = 12'b010001111011;
		if(({row_reg, col_reg}==18'b010100101010000010)) color_data = 12'b010101111011;
		if(({row_reg, col_reg}==18'b010100101010000011)) color_data = 12'b010101111010;
		if(({row_reg, col_reg}==18'b010100101010000100)) color_data = 12'b011001111000;
		if(({row_reg, col_reg}==18'b010100101010000101)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}==18'b010100101010000110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010100101010000111)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==18'b010100101010001000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100101010001001)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==18'b010100101010001010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100101010001011)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010100101010001100) && ({row_reg, col_reg}<18'b010100101010001110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010100101010001110) && ({row_reg, col_reg}<18'b010100101010010011)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010100101010010011) && ({row_reg, col_reg}<18'b010100101010100000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100101010100000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010100101010100001) && ({row_reg, col_reg}<18'b010100101010101001)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100101010101001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010100101010101010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010100101010101011) && ({row_reg, col_reg}<18'b010100101010101101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010100101010101101)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==18'b010100101010101110)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==18'b010100101010101111)) color_data = 12'b101010011000;
		if(({row_reg, col_reg}>=18'b010100101010110000) && ({row_reg, col_reg}<18'b010100101010110011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010100101010110011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010100101010110100)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010100101010110101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010100101010110110)) color_data = 12'b100110101001;
		if(({row_reg, col_reg}==18'b010100101010110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010100101010111000)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010100101010111001)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010100101010111010)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}>=18'b010100101010111011) && ({row_reg, col_reg}<18'b010100101011001011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100101011001011)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010100101011001100) && ({row_reg, col_reg}<18'b010100101011011110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010100101011011110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010100101011011111) && ({row_reg, col_reg}<18'b010100101011110010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010100101011110010) && ({row_reg, col_reg}<18'b010100101011110100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010100101011110100) && ({row_reg, col_reg}<18'b010100101011111000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100101011111000)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010100101011111001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010100101011111010) && ({row_reg, col_reg}<18'b010100101011111100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100101011111100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010100101011111101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010100101011111110)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}==18'b010100101011111111)) color_data = 12'b010101110110;
		if(({row_reg, col_reg}==18'b010100101100000000)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b010100101100000001)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}>=18'b010100101100000010) && ({row_reg, col_reg}<18'b010100101100000100)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010100101100000100)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010100101100000101)) color_data = 12'b011110111101;
		if(({row_reg, col_reg}==18'b010100101100000110)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b010100101100000111)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b010100101100001000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010100101100001001)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}>=18'b010100101100001010) && ({row_reg, col_reg}<18'b010100101100001100)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b010100101100001100)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}==18'b010100101100001101)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b010100101100001110)) color_data = 12'b011111001111;
		if(({row_reg, col_reg}==18'b010100101100001111)) color_data = 12'b011010111110;

		if(({row_reg, col_reg}>=18'b010100101100010000) && ({row_reg, col_reg}<18'b010100110000000000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010100110000000000) && ({row_reg, col_reg}<18'b010100110000000011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010100110000000011) && ({row_reg, col_reg}<18'b010100110000000110)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b010100110000000110) && ({row_reg, col_reg}<18'b010100110000001101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010100110000001101) && ({row_reg, col_reg}<18'b010100110000010000)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b010100110000010000) && ({row_reg, col_reg}<18'b010100110000010010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010100110000010010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b010100110000010011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010100110000010100) && ({row_reg, col_reg}<18'b010100110000010110)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}==18'b010100110000010110)) color_data = 12'b011111001110;
		if(({row_reg, col_reg}>=18'b010100110000010111) && ({row_reg, col_reg}<18'b010100110000011001)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010100110000011001)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}>=18'b010100110000011010) && ({row_reg, col_reg}<18'b010100110000011100)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010100110000011100) && ({row_reg, col_reg}<18'b010100110000100100)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010100110000100100)) color_data = 12'b100011111110;
		if(({row_reg, col_reg}==18'b010100110000100101)) color_data = 12'b100111111110;
		if(({row_reg, col_reg}==18'b010100110000100110)) color_data = 12'b100111101110;
		if(({row_reg, col_reg}==18'b010100110000100111)) color_data = 12'b100111101101;
		if(({row_reg, col_reg}==18'b010100110000101000)) color_data = 12'b101111101110;
		if(({row_reg, col_reg}==18'b010100110000101001)) color_data = 12'b100111001100;
		if(({row_reg, col_reg}==18'b010100110000101010)) color_data = 12'b010101110111;
		if(({row_reg, col_reg}>=18'b010100110000101011) && ({row_reg, col_reg}<18'b010100110000101101)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==18'b010100110000101101)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}>=18'b010100110000101110) && ({row_reg, col_reg}<18'b010100110000110000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010100110000110000)) color_data = 12'b011001110101;
		if(({row_reg, col_reg}==18'b010100110000110001)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}>=18'b010100110000110010) && ({row_reg, col_reg}<18'b010100110000110101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100110000110101)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==18'b010100110000110110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100110000110111)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010100110000111000) && ({row_reg, col_reg}<18'b010100110001000001)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010100110001000001) && ({row_reg, col_reg}<18'b010100110001000101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010100110001000101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010100110001000110) && ({row_reg, col_reg}<18'b010100110001001010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010100110001001010)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010100110001001011)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==18'b010100110001001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010100110001001101)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==18'b010100110001001110)) color_data = 12'b010101100111;
		if(({row_reg, col_reg}==18'b010100110001001111)) color_data = 12'b010001111000;
		if(({row_reg, col_reg}==18'b010100110001010000)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010100110001010001)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010100110001010010)) color_data = 12'b001101101101;
		if(({row_reg, col_reg}==18'b010100110001010011)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010100110001010100)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010100110001010101)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b010100110001010110) && ({row_reg, col_reg}<18'b010100110001011010)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010100110001011010)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010100110001011011)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b010100110001011100)) color_data = 12'b000101111011;
		if(({row_reg, col_reg}==18'b010100110001011101)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b010100110001011110)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010100110001011111)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}>=18'b010100110001100000) && ({row_reg, col_reg}<18'b010100110001100010)) color_data = 12'b101011101111;
		if(({row_reg, col_reg}==18'b010100110001100010)) color_data = 12'b100111011101;
		if(({row_reg, col_reg}==18'b010100110001100011)) color_data = 12'b100010111011;
		if(({row_reg, col_reg}==18'b010100110001100100)) color_data = 12'b100110111011;
		if(({row_reg, col_reg}==18'b010100110001100101)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b010100110001100110)) color_data = 12'b101010111011;
		if(({row_reg, col_reg}==18'b010100110001100111)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}==18'b010100110001101000)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==18'b010100110001101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010100110001101010) && ({row_reg, col_reg}<18'b010100110001101100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010100110001101100)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010100110001101101)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010100110001101110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010100110001101111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010100110001110000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010100110001110001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010100110001110010)) color_data = 12'b101010111010;
		if(({row_reg, col_reg}==18'b010100110001110011)) color_data = 12'b100110111011;
		if(({row_reg, col_reg}==18'b010100110001110100)) color_data = 12'b100110111100;
		if(({row_reg, col_reg}==18'b010100110001110101)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}==18'b010100110001110110)) color_data = 12'b010010001011;
		if(({row_reg, col_reg}==18'b010100110001110111)) color_data = 12'b001101111011;
		if(({row_reg, col_reg}==18'b010100110001111000)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b010100110001111001)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}==18'b010100110001111010)) color_data = 12'b001101111111;
		if(({row_reg, col_reg}==18'b010100110001111011)) color_data = 12'b001001111111;
		if(({row_reg, col_reg}==18'b010100110001111100)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b010100110001111101)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b010100110001111110) && ({row_reg, col_reg}<18'b010100110010000000)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010100110010000000)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010100110010000001)) color_data = 12'b010001111100;
		if(({row_reg, col_reg}==18'b010100110010000010)) color_data = 12'b010001111011;
		if(({row_reg, col_reg}==18'b010100110010000011)) color_data = 12'b010101111010;
		if(({row_reg, col_reg}==18'b010100110010000100)) color_data = 12'b010101111000;
		if(({row_reg, col_reg}==18'b010100110010000101)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==18'b010100110010000110)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}==18'b010100110010000111)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==18'b010100110010001000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010100110010001001)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==18'b010100110010001010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010100110010001011) && ({row_reg, col_reg}<18'b010100110010001111)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010100110010001111) && ({row_reg, col_reg}<18'b010100110010010010)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}==18'b010100110010010010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010100110010010011)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}>=18'b010100110010010100) && ({row_reg, col_reg}<18'b010100110010010110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010100110010010110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010100110010010111) && ({row_reg, col_reg}<18'b010100110010011011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010100110010011011) && ({row_reg, col_reg}<18'b010100110010011111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010100110010011111) && ({row_reg, col_reg}<18'b010100110010100001)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010100110010100001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010100110010100010) && ({row_reg, col_reg}<18'b010100110010100110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010100110010100110) && ({row_reg, col_reg}<18'b010100110010101001)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010100110010101001)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100110010101010)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010100110010101011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010100110010101100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010100110010101101)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==18'b010100110010101110)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==18'b010100110010101111)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}>=18'b010100110010110000) && ({row_reg, col_reg}<18'b010100110010110011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010100110010110011)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010100110010110100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010100110010110101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b010100110010110110) && ({row_reg, col_reg}<18'b010100110010111000)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010100110010111000)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b010100110010111001) && ({row_reg, col_reg}<18'b010100110010111100)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}>=18'b010100110010111100) && ({row_reg, col_reg}<18'b010100110011001011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100110011001011)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010100110011001100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010100110011001101)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b010100110011001110) && ({row_reg, col_reg}<18'b010100110011011111)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010100110011011111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010100110011100000) && ({row_reg, col_reg}<18'b010100110011110010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010100110011110010) && ({row_reg, col_reg}<18'b010100110011110100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010100110011110100) && ({row_reg, col_reg}<18'b010100110011111001)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100110011111001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010100110011111010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100110011111011)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010100110011111100) && ({row_reg, col_reg}<18'b010100110011111110)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}==18'b010100110011111110)) color_data = 12'b010101110110;
		if(({row_reg, col_reg}==18'b010100110011111111)) color_data = 12'b010001110110;
		if(({row_reg, col_reg}==18'b010100110100000000)) color_data = 12'b100011011110;
		if(({row_reg, col_reg}==18'b010100110100000001)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010100110100000010)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010100110100000011)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010100110100000100)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010100110100000101)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}==18'b010100110100000110)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}==18'b010100110100000111)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b010100110100001000)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}==18'b010100110100001001)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}==18'b010100110100001010)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010100110100001011)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b010100110100001100)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}==18'b010100110100001101)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b010100110100001110)) color_data = 12'b011111001110;
		if(({row_reg, col_reg}==18'b010100110100001111)) color_data = 12'b010110101101;
		if(({row_reg, col_reg}==18'b010100110100010000)) color_data = 12'b011010101110;

		if(({row_reg, col_reg}>=18'b010100110100010001) && ({row_reg, col_reg}<18'b010100111000000000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010100111000000000) && ({row_reg, col_reg}<18'b010100111000000010)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}>=18'b010100111000000010) && ({row_reg, col_reg}<18'b010100111000001001)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b010100111000001001) && ({row_reg, col_reg}<18'b010100111000001100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010100111000001100) && ({row_reg, col_reg}<18'b010100111000010000)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b010100111000010000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010100111000010001) && ({row_reg, col_reg}<18'b010100111000010011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010100111000010011)) color_data = 12'b011110111110;
		if(({row_reg, col_reg}==18'b010100111000010100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010100111000010101)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}==18'b010100111000010110)) color_data = 12'b011111001110;
		if(({row_reg, col_reg}>=18'b010100111000010111) && ({row_reg, col_reg}<18'b010100111000011001)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010100111000011001)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010100111000011010) && ({row_reg, col_reg}<18'b010100111000011100)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010100111000011100) && ({row_reg, col_reg}<18'b010100111000100011)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010100111000100011) && ({row_reg, col_reg}<18'b010100111000100111)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010100111000100111)) color_data = 12'b101011101111;
		if(({row_reg, col_reg}==18'b010100111000101000)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}==18'b010100111000101001)) color_data = 12'b100111001100;
		if(({row_reg, col_reg}==18'b010100111000101010)) color_data = 12'b010001110111;
		if(({row_reg, col_reg}==18'b010100111000101011)) color_data = 12'b010101111000;
		if(({row_reg, col_reg}==18'b010100111000101100)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==18'b010100111000101101)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}==18'b010100111000101110)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==18'b010100111000101111)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}>=18'b010100111000110000) && ({row_reg, col_reg}<18'b010100111000111010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100111000111010)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010100111000111011) && ({row_reg, col_reg}<18'b010100111001000110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100111001000110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010100111001000111) && ({row_reg, col_reg}<18'b010100111001001011)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}==18'b010100111001001011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010100111001001100)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==18'b010100111001001101)) color_data = 12'b010101100110;
		if(({row_reg, col_reg}==18'b010100111001001110)) color_data = 12'b010101111000;
		if(({row_reg, col_reg}==18'b010100111001001111)) color_data = 12'b010101111001;
		if(({row_reg, col_reg}==18'b010100111001010000)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010100111001010001)) color_data = 12'b010001111110;
		if(({row_reg, col_reg}>=18'b010100111001010010) && ({row_reg, col_reg}<18'b010100111001010100)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b010100111001010100) && ({row_reg, col_reg}<18'b010100111001010110)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010100111001010110)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b010100111001010111)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}==18'b010100111001011000)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b010100111001011001) && ({row_reg, col_reg}<18'b010100111001011100)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b010100111001011100)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b010100111001011101)) color_data = 12'b001110001011;
		if(({row_reg, col_reg}==18'b010100111001011110)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b010100111001011111)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}==18'b010100111001100000)) color_data = 12'b101011101111;
		if(({row_reg, col_reg}==18'b010100111001100001)) color_data = 12'b101111111111;
		if(({row_reg, col_reg}==18'b010100111001100010)) color_data = 12'b101011011101;
		if(({row_reg, col_reg}==18'b010100111001100011)) color_data = 12'b100010111011;
		if(({row_reg, col_reg}==18'b010100111001100100)) color_data = 12'b100110111011;
		if(({row_reg, col_reg}==18'b010100111001100101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010100111001100110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==18'b010100111001100111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010100111001101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010100111001101001)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010100111001101010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010100111001101011)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010100111001101100)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b010100111001101101) && ({row_reg, col_reg}<18'b010100111001101111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010100111001101111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010100111001110000)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010100111001110001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010100111001110010)) color_data = 12'b101010111010;
		if(({row_reg, col_reg}==18'b010100111001110011)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b010100111001110100)) color_data = 12'b100110111100;
		if(({row_reg, col_reg}==18'b010100111001110101)) color_data = 12'b011110011011;
		if(({row_reg, col_reg}==18'b010100111001110110)) color_data = 12'b010101111010;
		if(({row_reg, col_reg}==18'b010100111001110111)) color_data = 12'b010001111010;
		if(({row_reg, col_reg}==18'b010100111001111000)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}>=18'b010100111001111001) && ({row_reg, col_reg}<18'b010100111001111100)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b010100111001111100) && ({row_reg, col_reg}<18'b010100111010000000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010100111010000000) && ({row_reg, col_reg}<18'b010100111010000010)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010100111010000010)) color_data = 12'b001101111011;
		if(({row_reg, col_reg}==18'b010100111010000011)) color_data = 12'b001101111010;
		if(({row_reg, col_reg}==18'b010100111010000100)) color_data = 12'b010001101001;
		if(({row_reg, col_reg}==18'b010100111010000101)) color_data = 12'b010101111000;
		if(({row_reg, col_reg}==18'b010100111010000110)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==18'b010100111010000111)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}==18'b010100111010001000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010100111010001001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010100111010001010) && ({row_reg, col_reg}<18'b010100111010001111)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==18'b010100111010001111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010100111010010000) && ({row_reg, col_reg}<18'b010100111010010010)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==18'b010100111010010010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010100111010010011) && ({row_reg, col_reg}<18'b010100111010010101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100111010010101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010100111010010110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010100111010010111) && ({row_reg, col_reg}<18'b010100111010011001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010100111010011001) && ({row_reg, col_reg}<18'b010100111010011110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100111010011110)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==18'b010100111010011111)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}>=18'b010100111010100000) && ({row_reg, col_reg}<18'b010100111010100110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010100111010100110) && ({row_reg, col_reg}<18'b010100111010101000)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==18'b010100111010101000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010100111010101001) && ({row_reg, col_reg}<18'b010100111010101101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100111010101101)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==18'b010100111010101110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010100111010101111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010100111010110000) && ({row_reg, col_reg}<18'b010100111010110011)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}>=18'b010100111010110011) && ({row_reg, col_reg}<18'b010100111010110101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010100111010110101)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}>=18'b010100111010110110) && ({row_reg, col_reg}<18'b010100111010111000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010100111010111000)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b010100111010111001) && ({row_reg, col_reg}<18'b010100111010111100)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}>=18'b010100111010111100) && ({row_reg, col_reg}<18'b010100111011001011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100111011001011)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010100111011001100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010100111011001101) && ({row_reg, col_reg}<18'b010100111011001111)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b010100111011001111) && ({row_reg, col_reg}<18'b010100111011011110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010100111011011110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010100111011011111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010100111011100000) && ({row_reg, col_reg}<18'b010100111011111001)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010100111011111001)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010100111011111010) && ({row_reg, col_reg}<18'b010100111011111101)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}==18'b010100111011111101)) color_data = 12'b010101110110;
		if(({row_reg, col_reg}==18'b010100111011111110)) color_data = 12'b010001110110;
		if(({row_reg, col_reg}==18'b010100111011111111)) color_data = 12'b010010000111;
		if(({row_reg, col_reg}==18'b010100111100000000)) color_data = 12'b100011101110;
		if(({row_reg, col_reg}==18'b010100111100000001)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}==18'b010100111100000010)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010100111100000011)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010100111100000100)) color_data = 12'b100011101110;
		if(({row_reg, col_reg}==18'b010100111100000101)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}==18'b010100111100000110)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b010100111100000111)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b010100111100001000)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}==18'b010100111100001001)) color_data = 12'b011111001111;
		if(({row_reg, col_reg}>=18'b010100111100001010) && ({row_reg, col_reg}<18'b010100111100001100)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010100111100001100)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}==18'b010100111100001101)) color_data = 12'b101011101111;
		if(({row_reg, col_reg}==18'b010100111100001110)) color_data = 12'b011111001110;
		if(({row_reg, col_reg}==18'b010100111100001111)) color_data = 12'b010110101101;
		if(({row_reg, col_reg}==18'b010100111100010000)) color_data = 12'b011010101101;

		if(({row_reg, col_reg}>=18'b010100111100010001) && ({row_reg, col_reg}<18'b010101000000000001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010101000000000001) && ({row_reg, col_reg}<18'b010101000000000110)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b010101000000000110)) color_data = 12'b010110101111;
		if(({row_reg, col_reg}>=18'b010101000000000111) && ({row_reg, col_reg}<18'b010101000000001001)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b010101000000001001)) color_data = 12'b011010111111;
		if(({row_reg, col_reg}==18'b010101000000001010)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b010101000000001011) && ({row_reg, col_reg}<18'b010101000000010001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010101000000010001)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010101000000010010) && ({row_reg, col_reg}<18'b010101000000010101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010101000000010101)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==18'b010101000000010110)) color_data = 12'b011111001111;
		if(({row_reg, col_reg}>=18'b010101000000010111) && ({row_reg, col_reg}<18'b010101000000011001)) color_data = 12'b100011011111;
		if(({row_reg, col_reg}>=18'b010101000000011001) && ({row_reg, col_reg}<18'b010101000000011100)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}>=18'b010101000000011100) && ({row_reg, col_reg}<18'b010101000000100000)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010101000000100000) && ({row_reg, col_reg}<18'b010101000000100010)) color_data = 12'b011111101111;
		if(({row_reg, col_reg}==18'b010101000000100010)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010101000000100011)) color_data = 12'b011111101111;
		if(({row_reg, col_reg}==18'b010101000000100100)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}==18'b010101000000100101)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}>=18'b010101000000100110) && ({row_reg, col_reg}<18'b010101000000101001)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b010101000000101001)) color_data = 12'b011110111101;
		if(({row_reg, col_reg}==18'b010101000000101010)) color_data = 12'b001101111001;
		if(({row_reg, col_reg}>=18'b010101000000101011) && ({row_reg, col_reg}<18'b010101000000101101)) color_data = 12'b010101111001;
		if(({row_reg, col_reg}==18'b010101000000101101)) color_data = 12'b010101111000;
		if(({row_reg, col_reg}==18'b010101000000101110)) color_data = 12'b011001111000;
		if(({row_reg, col_reg}==18'b010101000000101111)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}>=18'b010101000000110000) && ({row_reg, col_reg}<18'b010101000001001000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010101000001001000)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==18'b010101000001001001)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010101000001001010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010101000001001011)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==18'b010101000001001100)) color_data = 12'b010101110111;
		if(({row_reg, col_reg}==18'b010101000001001101)) color_data = 12'b010001110111;
		if(({row_reg, col_reg}==18'b010101000001001110)) color_data = 12'b010110001001;
		if(({row_reg, col_reg}==18'b010101000001001111)) color_data = 12'b010010001001;
		if(({row_reg, col_reg}==18'b010101000001010000)) color_data = 12'b001001101100;
		if(({row_reg, col_reg}==18'b010101000001010001)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b010101000001010010) && ({row_reg, col_reg}<18'b010101000001010100)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}>=18'b010101000001010100) && ({row_reg, col_reg}<18'b010101000001011000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010101000001011000)) color_data = 12'b001001101101;
		if(({row_reg, col_reg}>=18'b010101000001011001) && ({row_reg, col_reg}<18'b010101000001011011)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010101000001011011)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010101000001011100)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010101000001011101)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b010101000001011110)) color_data = 12'b100111011111;
		if(({row_reg, col_reg}==18'b010101000001011111)) color_data = 12'b101011101111;
		if(({row_reg, col_reg}==18'b010101000001100000)) color_data = 12'b101011011110;
		if(({row_reg, col_reg}==18'b010101000001100001)) color_data = 12'b101111101111;
		if(({row_reg, col_reg}==18'b010101000001100010)) color_data = 12'b101111011101;
		if(({row_reg, col_reg}==18'b010101000001100011)) color_data = 12'b100110111011;
		if(({row_reg, col_reg}>=18'b010101000001100100) && ({row_reg, col_reg}<18'b010101000001100110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010101000001100110)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==18'b010101000001100111)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==18'b010101000001101000)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010101000001101001) && ({row_reg, col_reg}<18'b010101000001101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010101000001101100)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}>=18'b010101000001101101) && ({row_reg, col_reg}<18'b010101000001110000)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010101000001110000)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b010101000001110001) && ({row_reg, col_reg}<18'b010101000001110011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010101000001110011)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b010101000001110100)) color_data = 12'b101010111100;
		if(({row_reg, col_reg}==18'b010101000001110101)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}==18'b010101000001110110)) color_data = 12'b011010001010;
		if(({row_reg, col_reg}==18'b010101000001110111)) color_data = 12'b010101111010;
		if(({row_reg, col_reg}>=18'b010101000001111000) && ({row_reg, col_reg}<18'b010101000001111010)) color_data = 12'b010001111011;
		if(({row_reg, col_reg}==18'b010101000001111010)) color_data = 12'b010001111100;
		if(({row_reg, col_reg}>=18'b010101000001111011) && ({row_reg, col_reg}<18'b010101000010000000)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b010101000010000000)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}>=18'b010101000010000001) && ({row_reg, col_reg}<18'b010101000010000011)) color_data = 12'b001110001011;
		if(({row_reg, col_reg}==18'b010101000010000011)) color_data = 12'b010110011100;
		if(({row_reg, col_reg}==18'b010101000010000100)) color_data = 12'b010001111010;
		if(({row_reg, col_reg}==18'b010101000010000101)) color_data = 12'b010001111001;
		if(({row_reg, col_reg}==18'b010101000010000110)) color_data = 12'b010101111001;
		if(({row_reg, col_reg}==18'b010101000010000111)) color_data = 12'b011001111000;
		if(({row_reg, col_reg}==18'b010101000010001000)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}>=18'b010101000010001001) && ({row_reg, col_reg}<18'b010101000010001011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010101000010001011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010101000010001100)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010101000010001101) && ({row_reg, col_reg}<18'b010101000010011110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010101000010011110) && ({row_reg, col_reg}<18'b010101000010100000)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}>=18'b010101000010100000) && ({row_reg, col_reg}<18'b010101000010100010)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010101000010100010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010101000010100011) && ({row_reg, col_reg}<18'b010101000010100101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010101000010100101) && ({row_reg, col_reg}<18'b010101000010101000)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010101000010101000)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==18'b010101000010101001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010101000010101010)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==18'b010101000010101011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010101000010101100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010101000010101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010101000010101110)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==18'b010101000010101111)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}>=18'b010101000010110000) && ({row_reg, col_reg}<18'b010101000010110100)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==18'b010101000010110100)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}==18'b010101000010110101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010101000010110110)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==18'b010101000010110111)) color_data = 12'b100110001001;
		if(({row_reg, col_reg}>=18'b010101000010111000) && ({row_reg, col_reg}<18'b010101000010111010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010101000010111010)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010101000010111011)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}>=18'b010101000010111100) && ({row_reg, col_reg}<18'b010101000010111110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010101000010111110) && ({row_reg, col_reg}<18'b010101000011000000)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010101000011000000) && ({row_reg, col_reg}<18'b010101000011001011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010101000011001011)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010101000011001100) && ({row_reg, col_reg}<18'b010101000011011000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010101000011011000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010101000011011001) && ({row_reg, col_reg}<18'b010101000011011110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010101000011011110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010101000011011111) && ({row_reg, col_reg}<18'b010101000011110000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010101000011110000)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}>=18'b010101000011110001) && ({row_reg, col_reg}<18'b010101000011111000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010101000011111000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010101000011111001)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010101000011111010)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}==18'b010101000011111011)) color_data = 12'b010101100110;
		if(({row_reg, col_reg}==18'b010101000011111100)) color_data = 12'b011010000111;
		if(({row_reg, col_reg}==18'b010101000011111101)) color_data = 12'b010001110111;
		if(({row_reg, col_reg}==18'b010101000011111110)) color_data = 12'b010010000111;
		if(({row_reg, col_reg}==18'b010101000011111111)) color_data = 12'b010010011000;
		if(({row_reg, col_reg}==18'b010101000100000000)) color_data = 12'b011111011110;
		if(({row_reg, col_reg}==18'b010101000100000001)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010101000100000010)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010101000100000011)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010101000100000100)) color_data = 12'b100011101110;
		if(({row_reg, col_reg}==18'b010101000100000101)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}==18'b010101000100000110)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b010101000100000111)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b010101000100001000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010101000100001001)) color_data = 12'b011111001111;
		if(({row_reg, col_reg}>=18'b010101000100001010) && ({row_reg, col_reg}<18'b010101000100001110)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b010101000100001110)) color_data = 12'b011111001110;
		if(({row_reg, col_reg}==18'b010101000100001111)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}>=18'b010101000100010000) && ({row_reg, col_reg}<18'b010101000100010010)) color_data = 12'b011010101110;

		if(({row_reg, col_reg}==18'b010101000100010010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010101001000000000) && ({row_reg, col_reg}<18'b010101001000000011)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b010101001000000011)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b010101001000000100) && ({row_reg, col_reg}<18'b010101001000000110)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b010101001000000110)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010101001000000111)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b010101001000001000)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==18'b010101001000001001)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b010101001000001010) && ({row_reg, col_reg}<18'b010101001000001111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010101001000001111) && ({row_reg, col_reg}<18'b010101001000010010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010101001000010010) && ({row_reg, col_reg}<18'b010101001000010110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010101001000010110)) color_data = 12'b010110101101;
		if(({row_reg, col_reg}>=18'b010101001000010111) && ({row_reg, col_reg}<18'b010101001000011001)) color_data = 12'b010010011101;
		if(({row_reg, col_reg}==18'b010101001000011001)) color_data = 12'b001110011100;
		if(({row_reg, col_reg}==18'b010101001000011010)) color_data = 12'b001110011011;
		if(({row_reg, col_reg}==18'b010101001000011011)) color_data = 12'b011111011110;
		if(({row_reg, col_reg}==18'b010101001000011100)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010101001000011101)) color_data = 12'b100011111110;
		if(({row_reg, col_reg}>=18'b010101001000011110) && ({row_reg, col_reg}<18'b010101001000100000)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010101001000100000)) color_data = 12'b010010101100;
		if(({row_reg, col_reg}==18'b010101001000100001)) color_data = 12'b001010011011;
		if(({row_reg, col_reg}==18'b010101001000100010)) color_data = 12'b001110011100;
		if(({row_reg, col_reg}>=18'b010101001000100011) && ({row_reg, col_reg}<18'b010101001000100110)) color_data = 12'b001110011101;
		if(({row_reg, col_reg}>=18'b010101001000100110) && ({row_reg, col_reg}<18'b010101001000101000)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b010101001000101000)) color_data = 12'b010010011101;
		if(({row_reg, col_reg}==18'b010101001000101001)) color_data = 12'b010010001100;
		if(({row_reg, col_reg}==18'b010101001000101010)) color_data = 12'b001101111011;
		if(({row_reg, col_reg}==18'b010101001000101011)) color_data = 12'b010010001011;
		if(({row_reg, col_reg}==18'b010101001000101100)) color_data = 12'b010001111010;
		if(({row_reg, col_reg}==18'b010101001000101101)) color_data = 12'b010101111001;
		if(({row_reg, col_reg}==18'b010101001000101110)) color_data = 12'b011001101001;
		if(({row_reg, col_reg}==18'b010101001000101111)) color_data = 12'b011001101000;
		if(({row_reg, col_reg}==18'b010101001000110000)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010101001000110001) && ({row_reg, col_reg}<18'b010101001000110110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010101001000110110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010101001000110111) && ({row_reg, col_reg}<18'b010101001000111001)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}>=18'b010101001000111001) && ({row_reg, col_reg}<18'b010101001001001010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010101001001001010)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==18'b010101001001001011)) color_data = 12'b101011001100;
		if(({row_reg, col_reg}==18'b010101001001001100)) color_data = 12'b101011011101;
		if(({row_reg, col_reg}==18'b010101001001001101)) color_data = 12'b100111011101;
		if(({row_reg, col_reg}==18'b010101001001001110)) color_data = 12'b100111011110;
		if(({row_reg, col_reg}==18'b010101001001001111)) color_data = 12'b011110111101;
		if(({row_reg, col_reg}==18'b010101001001010000)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b010101001001010001)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b010101001001010010) && ({row_reg, col_reg}<18'b010101001001010110)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010101001001010110)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010101001001010111)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010101001001011000)) color_data = 12'b001101111111;
		if(({row_reg, col_reg}==18'b010101001001011001)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b010101001001011010)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010101001001011011)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010101001001011100)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010101001001011101)) color_data = 12'b010010001011;
		if(({row_reg, col_reg}==18'b010101001001011110)) color_data = 12'b011110111101;
		if(({row_reg, col_reg}==18'b010101001001011111)) color_data = 12'b100010111101;
		if(({row_reg, col_reg}>=18'b010101001001100000) && ({row_reg, col_reg}<18'b010101001001100010)) color_data = 12'b100110111011;
		if(({row_reg, col_reg}==18'b010101001001100010)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}>=18'b010101001001100011) && ({row_reg, col_reg}<18'b010101001001100110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010101001001100110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010101001001100111)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}>=18'b010101001001101000) && ({row_reg, col_reg}<18'b010101001001101010)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010101001001101010)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}==18'b010101001001101011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010101001001101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010101001001101101)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b010101001001101110) && ({row_reg, col_reg}<18'b010101001001110000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010101001001110000)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010101001001110001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010101001001110010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010101001001110011)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}==18'b010101001001110100)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}>=18'b010101001001110101) && ({row_reg, col_reg}<18'b010101001001110111)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b010101001001110111)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b010101001001111000)) color_data = 12'b100010111100;
		if(({row_reg, col_reg}==18'b010101001001111001)) color_data = 12'b100010111101;
		if(({row_reg, col_reg}==18'b010101001001111010)) color_data = 12'b100011001110;
		if(({row_reg, col_reg}==18'b010101001001111011)) color_data = 12'b100111011111;
		if(({row_reg, col_reg}==18'b010101001001111100)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}>=18'b010101001001111101) && ({row_reg, col_reg}<18'b010101001010000000)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010101001010000000)) color_data = 12'b011111101111;
		if(({row_reg, col_reg}>=18'b010101001010000001) && ({row_reg, col_reg}<18'b010101001010000011)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010101001010000011)) color_data = 12'b100011011111;
		if(({row_reg, col_reg}==18'b010101001010000100)) color_data = 12'b010110011100;
		if(({row_reg, col_reg}==18'b010101001010000101)) color_data = 12'b001101111011;
		if(({row_reg, col_reg}==18'b010101001010000110)) color_data = 12'b010001111011;
		if(({row_reg, col_reg}==18'b010101001010000111)) color_data = 12'b010101111010;
		if(({row_reg, col_reg}==18'b010101001010001000)) color_data = 12'b011001111000;
		if(({row_reg, col_reg}==18'b010101001010001001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010101001010001010)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010101001010001011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010101001010001100) && ({row_reg, col_reg}<18'b010101001010010010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010101001010010010)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}>=18'b010101001010010011) && ({row_reg, col_reg}<18'b010101001010100000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010101001010100000)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==18'b010101001010100001)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}>=18'b010101001010100010) && ({row_reg, col_reg}<18'b010101001010100111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010101001010100111)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==18'b010101001010101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010101001010101001) && ({row_reg, col_reg}<18'b010101001010101011)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==18'b010101001010101011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010101001010101100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010101001010101101)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}==18'b010101001010101110)) color_data = 12'b100010011011;
		if(({row_reg, col_reg}==18'b010101001010101111)) color_data = 12'b011110001010;
		if(({row_reg, col_reg}==18'b010101001010110000)) color_data = 12'b011001111100;
		if(({row_reg, col_reg}==18'b010101001010110001)) color_data = 12'b010101111011;
		if(({row_reg, col_reg}==18'b010101001010110010)) color_data = 12'b011001111011;
		if(({row_reg, col_reg}==18'b010101001010110011)) color_data = 12'b011101111010;
		if(({row_reg, col_reg}==18'b010101001010110100)) color_data = 12'b011101111001;
		if(({row_reg, col_reg}==18'b010101001010110101)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==18'b010101001010110110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010101001010110111) && ({row_reg, col_reg}<18'b010101001010111001)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010101001010111001) && ({row_reg, col_reg}<18'b010101001010111110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010101001010111110) && ({row_reg, col_reg}<18'b010101001011000000)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010101001011000000) && ({row_reg, col_reg}<18'b010101001011001100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010101001011001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010101001011001101)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010101001011001110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010101001011001111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010101001011010000) && ({row_reg, col_reg}<18'b010101001011010101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010101001011010101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010101001011010110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010101001011010111) && ({row_reg, col_reg}<18'b010101001011011001)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010101001011011001)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010101001011011010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010101001011011011) && ({row_reg, col_reg}<18'b010101001011011110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010101001011011110) && ({row_reg, col_reg}<18'b010101001011110110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010101001011110110) && ({row_reg, col_reg}<18'b010101001011111001)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010101001011111001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010101001011111010)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==18'b010101001011111011)) color_data = 12'b100110111011;
		if(({row_reg, col_reg}==18'b010101001011111100)) color_data = 12'b101111101110;
		if(({row_reg, col_reg}>=18'b010101001011111101) && ({row_reg, col_reg}<18'b010101001011111111)) color_data = 12'b100111011101;
		if(({row_reg, col_reg}==18'b010101001011111111)) color_data = 12'b100011011100;
		if(({row_reg, col_reg}>=18'b010101001100000000) && ({row_reg, col_reg}<18'b010101001100000011)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010101001100000011)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010101001100000100)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010101001100000101)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}==18'b010101001100000110)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}==18'b010101001100000111)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b010101001100001000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010101001100001001)) color_data = 12'b011110111110;
		if(({row_reg, col_reg}==18'b010101001100001010)) color_data = 12'b011111001111;
		if(({row_reg, col_reg}==18'b010101001100001011)) color_data = 12'b011110111110;
		if(({row_reg, col_reg}==18'b010101001100001100)) color_data = 12'b011111001110;
		if(({row_reg, col_reg}==18'b010101001100001101)) color_data = 12'b011110111110;
		if(({row_reg, col_reg}==18'b010101001100001110)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}==18'b010101001100001111)) color_data = 12'b011010101101;

		if(({row_reg, col_reg}>=18'b010101001100010000) && ({row_reg, col_reg}<18'b010101010000000000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010101010000000000) && ({row_reg, col_reg}<18'b010101010000000100)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010101010000000100)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010101010000000101)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010101010000000110)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010101010000000111)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010101010000001000)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==18'b010101010000001001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010101010000001010)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}>=18'b010101010000001011) && ({row_reg, col_reg}<18'b010101010000001111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010101010000001111)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}==18'b010101010000010000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010101010000010001) && ({row_reg, col_reg}<18'b010101010000010011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010101010000010011) && ({row_reg, col_reg}<18'b010101010000010110)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b010101010000010110)) color_data = 12'b010110011101;
		if(({row_reg, col_reg}>=18'b010101010000010111) && ({row_reg, col_reg}<18'b010101010000011010)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010101010000011010)) color_data = 12'b001001111010;
		if(({row_reg, col_reg}==18'b010101010000011011)) color_data = 12'b011011001101;
		if(({row_reg, col_reg}==18'b010101010000011100)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010101010000011101)) color_data = 12'b100011111110;
		if(({row_reg, col_reg}==18'b010101010000011110)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010101010000011111)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010101010000100000)) color_data = 12'b001110011100;
		if(({row_reg, col_reg}==18'b010101010000100001)) color_data = 12'b000101111010;
		if(({row_reg, col_reg}==18'b010101010000100010)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}>=18'b010101010000100011) && ({row_reg, col_reg}<18'b010101010000100101)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b010101010000100101) && ({row_reg, col_reg}<18'b010101010000100111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010101010000100111)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b010101010000101000) && ({row_reg, col_reg}<18'b010101010000101010)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010101010000101010)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b010101010000101011)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b010101010000101100)) color_data = 12'b001101111011;
		if(({row_reg, col_reg}==18'b010101010000101101)) color_data = 12'b010001111010;
		if(({row_reg, col_reg}==18'b010101010000101110)) color_data = 12'b010101101001;
		if(({row_reg, col_reg}==18'b010101010000101111)) color_data = 12'b011001101001;
		if(({row_reg, col_reg}>=18'b010101010000110000) && ({row_reg, col_reg}<18'b010101010000110010)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010101010000110010) && ({row_reg, col_reg}<18'b010101010000110100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010101010000110100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010101010000110101)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==18'b010101010000110110)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}==18'b010101010000110111)) color_data = 12'b011001110101;
		if(({row_reg, col_reg}==18'b010101010000111000)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}==18'b010101010000111001)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}>=18'b010101010000111010) && ({row_reg, col_reg}<18'b010101010001001001)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010101010001001001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010101010001001010)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==18'b010101010001001011)) color_data = 12'b101111011101;
		if(({row_reg, col_reg}==18'b010101010001001100)) color_data = 12'b101111111111;
		if(({row_reg, col_reg}==18'b010101010001001101)) color_data = 12'b101011101110;
		if(({row_reg, col_reg}==18'b010101010001001110)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}==18'b010101010001001111)) color_data = 12'b100011001110;
		if(({row_reg, col_reg}==18'b010101010001010000)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b010101010001010001)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}>=18'b010101010001010010) && ({row_reg, col_reg}<18'b010101010001010101)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010101010001010101) && ({row_reg, col_reg}<18'b010101010001011000)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010101010001011000)) color_data = 12'b001001111111;
		if(({row_reg, col_reg}==18'b010101010001011001)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b010101010001011010)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010101010001011011)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010101010001011100)) color_data = 12'b001110001011;
		if(({row_reg, col_reg}==18'b010101010001011101)) color_data = 12'b010001111011;
		if(({row_reg, col_reg}==18'b010101010001011110)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}==18'b010101010001011111)) color_data = 12'b100110111100;
		if(({row_reg, col_reg}==18'b010101010001100000)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b010101010001100001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010101010001100010)) color_data = 12'b101010111011;
		if(({row_reg, col_reg}==18'b010101010001100011)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}>=18'b010101010001100100) && ({row_reg, col_reg}<18'b010101010001100111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010101010001100111)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010101010001101000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010101010001101001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010101010001101010)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010101010001101011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010101010001101100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010101010001101101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010101010001101110) && ({row_reg, col_reg}<18'b010101010001110000)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==18'b010101010001110000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010101010001110001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010101010001110010)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}>=18'b010101010001110011) && ({row_reg, col_reg}<18'b010101010001110101)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}==18'b010101010001110101)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==18'b010101010001110110)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b010101010001110111)) color_data = 12'b101010111011;
		if(({row_reg, col_reg}>=18'b010101010001111000) && ({row_reg, col_reg}<18'b010101010001111010)) color_data = 12'b100110111011;
		if(({row_reg, col_reg}==18'b010101010001111010)) color_data = 12'b100111001100;
		if(({row_reg, col_reg}==18'b010101010001111011)) color_data = 12'b101011101110;
		if(({row_reg, col_reg}==18'b010101010001111100)) color_data = 12'b101011111110;
		if(({row_reg, col_reg}>=18'b010101010001111101) && ({row_reg, col_reg}<18'b010101010001111111)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010101010001111111) && ({row_reg, col_reg}<18'b010101010010000100)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010101010010000100)) color_data = 12'b010110101101;
		if(({row_reg, col_reg}==18'b010101010010000101)) color_data = 12'b001101101100;
		if(({row_reg, col_reg}==18'b010101010010000110)) color_data = 12'b010001101100;
		if(({row_reg, col_reg}==18'b010101010010000111)) color_data = 12'b010101101011;
		if(({row_reg, col_reg}==18'b010101010010001000)) color_data = 12'b010101101001;
		if(({row_reg, col_reg}==18'b010101010010001001)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==18'b010101010010001010)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}==18'b010101010010001011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010101010010001100) && ({row_reg, col_reg}<18'b010101010010001111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010101010010001111)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}>=18'b010101010010010000) && ({row_reg, col_reg}<18'b010101010010100000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010101010010100000)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010101010010100001)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010101010010100010) && ({row_reg, col_reg}<18'b010101010010100111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b010101010010100111) && ({row_reg, col_reg}<18'b010101010010101011)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==18'b010101010010101011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010101010010101100)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==18'b010101010010101101)) color_data = 12'b101110111100;
		if(({row_reg, col_reg}==18'b010101010010101110)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==18'b010101010010101111)) color_data = 12'b010101111010;
		if(({row_reg, col_reg}==18'b010101010010110000)) color_data = 12'b010001101100;
		if(({row_reg, col_reg}==18'b010101010010110001)) color_data = 12'b010001101011;
		if(({row_reg, col_reg}==18'b010101010010110010)) color_data = 12'b010101101011;
		if(({row_reg, col_reg}==18'b010101010010110011)) color_data = 12'b010101101010;
		if(({row_reg, col_reg}==18'b010101010010110100)) color_data = 12'b010101101000;
		if(({row_reg, col_reg}>=18'b010101010010110101) && ({row_reg, col_reg}<18'b010101010010110111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010101010010110111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010101010010111000) && ({row_reg, col_reg}<18'b010101010010111010)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010101010010111010) && ({row_reg, col_reg}<18'b010101010011010000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010101010011010000) && ({row_reg, col_reg}<18'b010101010011010101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010101010011010101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010101010011010110) && ({row_reg, col_reg}<18'b010101010011110011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010101010011110011)) color_data = 12'b100001100110;
		if(({row_reg, col_reg}>=18'b010101010011110100) && ({row_reg, col_reg}<18'b010101010011110110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010101010011110110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010101010011110111) && ({row_reg, col_reg}<18'b010101010011111001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010101010011111001)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}==18'b010101010011111010)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==18'b010101010011111011)) color_data = 12'b100110111100;
		if(({row_reg, col_reg}==18'b010101010011111100)) color_data = 12'b101111111111;
		if(({row_reg, col_reg}>=18'b010101010011111101) && ({row_reg, col_reg}<18'b010101010011111111)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}==18'b010101010011111111)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010101010100000000) && ({row_reg, col_reg}<18'b010101010100000010)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010101010100000010) && ({row_reg, col_reg}<18'b010101010100000100)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010101010100000100)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010101010100000101)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}==18'b010101010100000110)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}==18'b010101010100000111)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b010101010100001000)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}==18'b010101010100001001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010101010100001010) && ({row_reg, col_reg}<18'b010101010100010000)) color_data = 12'b011010101101;

		if(({row_reg, col_reg}>=18'b010101010100010000) && ({row_reg, col_reg}<18'b010101011000000000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010101011000000000) && ({row_reg, col_reg}<18'b010101011000000010)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010101011000000010)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b010101011000000011)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010101011000000100)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b010101011000000101)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010101011000000110)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010101011000000111)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b010101011000001000)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==18'b010101011000001001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010101011000001010)) color_data = 12'b011110111111;
		if(({row_reg, col_reg}==18'b010101011000001011)) color_data = 12'b011110111110;
		if(({row_reg, col_reg}==18'b010101011000001100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010101011000001101) && ({row_reg, col_reg}<18'b010101011000010000)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}>=18'b010101011000010000) && ({row_reg, col_reg}<18'b010101011000010100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010101011000010100) && ({row_reg, col_reg}<18'b010101011000010110)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b010101011000010110)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==18'b010101011000010111)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010101011000011000)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010101011000011001)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010101011000011010)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b010101011000011011)) color_data = 12'b011011001110;
		if(({row_reg, col_reg}>=18'b010101011000011100) && ({row_reg, col_reg}<18'b010101011000100000)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010101011000100000)) color_data = 12'b001110011100;
		if(({row_reg, col_reg}==18'b010101011000100001)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b010101011000100010)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}>=18'b010101011000100011) && ({row_reg, col_reg}<18'b010101011000100101)) color_data = 12'b001010001101;
		if(({row_reg, col_reg}>=18'b010101011000100101) && ({row_reg, col_reg}<18'b010101011000100111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010101011000100111) && ({row_reg, col_reg}<18'b010101011000101001)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010101011000101001)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010101011000101010)) color_data = 12'b001010001101;
		if(({row_reg, col_reg}==18'b010101011000101011)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b010101011000101100)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b010101011000101101)) color_data = 12'b010001111011;
		if(({row_reg, col_reg}==18'b010101011000101110)) color_data = 12'b010101111010;
		if(({row_reg, col_reg}==18'b010101011000101111)) color_data = 12'b010101111001;
		if(({row_reg, col_reg}>=18'b010101011000110000) && ({row_reg, col_reg}<18'b010101011000110011)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}==18'b010101011000110011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010101011000110100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010101011000110101) && ({row_reg, col_reg}<18'b010101011000110111)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}==18'b010101011000110111)) color_data = 12'b010101100110;
		if(({row_reg, col_reg}>=18'b010101011000111000) && ({row_reg, col_reg}<18'b010101011000111010)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}>=18'b010101011000111010) && ({row_reg, col_reg}<18'b010101011000111100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010101011000111100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010101011000111101)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010101011000111110) && ({row_reg, col_reg}<18'b010101011001000000)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}==18'b010101011001000000)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==18'b010101011001000001)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}==18'b010101011001000010)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==18'b010101011001000011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010101011001000100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010101011001000101) && ({row_reg, col_reg}<18'b010101011001000111)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}>=18'b010101011001000111) && ({row_reg, col_reg}<18'b010101011001001001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010101011001001001)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==18'b010101011001001010)) color_data = 12'b011001111000;
		if(({row_reg, col_reg}==18'b010101011001001011)) color_data = 12'b101011011101;
		if(({row_reg, col_reg}==18'b010101011001001100)) color_data = 12'b101011111110;
		if(({row_reg, col_reg}==18'b010101011001001101)) color_data = 12'b100111101110;
		if(({row_reg, col_reg}==18'b010101011001001110)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}==18'b010101011001001111)) color_data = 12'b011111001110;
		if(({row_reg, col_reg}==18'b010101011001010000)) color_data = 12'b000101111010;
		if(({row_reg, col_reg}==18'b010101011001010001)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b010101011001010010)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b010101011001010011)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}>=18'b010101011001010100) && ({row_reg, col_reg}<18'b010101011001010110)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010101011001010110) && ({row_reg, col_reg}<18'b010101011001011000)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010101011001011000)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b010101011001011001)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010101011001011010)) color_data = 12'b001010001101;
		if(({row_reg, col_reg}==18'b010101011001011011)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b010101011001011100)) color_data = 12'b001101111010;
		if(({row_reg, col_reg}==18'b010101011001011101)) color_data = 12'b010010001010;
		if(({row_reg, col_reg}==18'b010101011001011110)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b010101011001011111)) color_data = 12'b100110111100;
		if(({row_reg, col_reg}>=18'b010101011001100000) && ({row_reg, col_reg}<18'b010101011001100010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010101011001100010)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==18'b010101011001100011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010101011001100100)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}>=18'b010101011001100101) && ({row_reg, col_reg}<18'b010101011001100111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010101011001100111)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==18'b010101011001101000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010101011001101001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010101011001101010)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010101011001101011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010101011001101100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010101011001101101)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b010101011001101110) && ({row_reg, col_reg}<18'b010101011001110000)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==18'b010101011001110000)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010101011001110001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010101011001110010)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010101011001110011) && ({row_reg, col_reg}<18'b010101011001110110)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==18'b010101011001110110)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b010101011001110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010101011001111000)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==18'b010101011001111001)) color_data = 12'b100110111010;
		if(({row_reg, col_reg}==18'b010101011001111010)) color_data = 12'b100111001011;
		if(({row_reg, col_reg}==18'b010101011001111011)) color_data = 12'b101111101101;
		if(({row_reg, col_reg}==18'b010101011001111100)) color_data = 12'b101011101101;
		if(({row_reg, col_reg}==18'b010101011001111101)) color_data = 12'b100111111110;
		if(({row_reg, col_reg}==18'b010101011001111110)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010101011001111111) && ({row_reg, col_reg}<18'b010101011010000100)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010101011010000100)) color_data = 12'b010010011101;
		if(({row_reg, col_reg}==18'b010101011010000101)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010101011010000110)) color_data = 12'b010001111110;
		if(({row_reg, col_reg}==18'b010101011010000111)) color_data = 12'b010001111100;
		if(({row_reg, col_reg}==18'b010101011010001000)) color_data = 12'b010101111010;
		if(({row_reg, col_reg}==18'b010101011010001001)) color_data = 12'b010101101000;
		if(({row_reg, col_reg}>=18'b010101011010001010) && ({row_reg, col_reg}<18'b010101011010001100)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==18'b010101011010001100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010101011010001101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010101011010001110)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}==18'b010101011010001111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010101011010010000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010101011010010001)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010101011010010010) && ({row_reg, col_reg}<18'b010101011010010101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010101011010010101) && ({row_reg, col_reg}<18'b010101011010010111)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==18'b010101011010010111)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}>=18'b010101011010011000) && ({row_reg, col_reg}<18'b010101011010011100)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010101011010011100) && ({row_reg, col_reg}<18'b010101011010011110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010101011010011110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010101011010011111)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==18'b010101011010100000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010101011010100001) && ({row_reg, col_reg}<18'b010101011010100100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010101011010100100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010101011010100101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010101011010100110)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b010101011010100111)) color_data = 12'b101010111011;
		if(({row_reg, col_reg}==18'b010101011010101000)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b010101011010101001)) color_data = 12'b101110101100;
		if(({row_reg, col_reg}==18'b010101011010101010)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b010101011010101011)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==18'b010101011010101100)) color_data = 12'b101010101011;
		if(({row_reg, col_reg}==18'b010101011010101101)) color_data = 12'b101010111100;
		if(({row_reg, col_reg}==18'b010101011010101110)) color_data = 12'b100010101101;
		if(({row_reg, col_reg}==18'b010101011010101111)) color_data = 12'b010101111010;
		if(({row_reg, col_reg}==18'b010101011010110000)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}>=18'b010101011010110001) && ({row_reg, col_reg}<18'b010101011010110011)) color_data = 12'b010001111100;
		if(({row_reg, col_reg}==18'b010101011010110011)) color_data = 12'b010101111010;
		if(({row_reg, col_reg}==18'b010101011010110100)) color_data = 12'b010101111000;
		if(({row_reg, col_reg}>=18'b010101011010110101) && ({row_reg, col_reg}<18'b010101011010110111)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==18'b010101011010110111)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}>=18'b010101011010111000) && ({row_reg, col_reg}<18'b010101011010111011)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010101011010111011) && ({row_reg, col_reg}<18'b010101011010111110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010101011010111110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010101011010111111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010101011011000000) && ({row_reg, col_reg}<18'b010101011011010000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010101011011010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010101011011010001) && ({row_reg, col_reg}<18'b010101011011010101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010101011011010101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010101011011010110) && ({row_reg, col_reg}<18'b010101011011101011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010101011011101011)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010101011011101100) && ({row_reg, col_reg}<18'b010101011011110010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010101011011110010) && ({row_reg, col_reg}<18'b010101011011110100)) color_data = 12'b100001100110;
		if(({row_reg, col_reg}==18'b010101011011110100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010101011011110101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010101011011110110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010101011011110111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010101011011111000)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}==18'b010101011011111001)) color_data = 12'b011110001000;
		if(({row_reg, col_reg}==18'b010101011011111010)) color_data = 12'b010001100111;
		if(({row_reg, col_reg}==18'b010101011011111011)) color_data = 12'b100010111100;
		if(({row_reg, col_reg}==18'b010101011011111100)) color_data = 12'b101111111111;
		if(({row_reg, col_reg}==18'b010101011011111101)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b010101011011111110)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010101011011111111)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}>=18'b010101011100000000) && ({row_reg, col_reg}<18'b010101011100000010)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010101011100000010) && ({row_reg, col_reg}<18'b010101011100000100)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010101011100000100)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010101011100000101)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}==18'b010101011100000110)) color_data = 12'b010110101101;
		if(({row_reg, col_reg}==18'b010101011100000111)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}>=18'b010101011100001000) && ({row_reg, col_reg}<18'b010101011100001011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010101011100001011)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}>=18'b010101011100001100) && ({row_reg, col_reg}<18'b010101011100001111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010101011100001111)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b010101011100010000) && ({row_reg, col_reg}<18'b010101100000000000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010101100000000000)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010101100000000001)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010101100000000010)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010101100000000011)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b010101100000000100) && ({row_reg, col_reg}<18'b010101100000000111)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010101100000000111)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b010101100000001000)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}>=18'b010101100000001001) && ({row_reg, col_reg}<18'b010101100000001111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010101100000001111)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b010101100000010000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010101100000010001)) color_data = 12'b011110111110;
		if(({row_reg, col_reg}>=18'b010101100000010010) && ({row_reg, col_reg}<18'b010101100000010100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010101100000010100)) color_data = 12'b011110111111;
		if(({row_reg, col_reg}==18'b010101100000010101)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b010101100000010110)) color_data = 12'b010010011110;
		if(({row_reg, col_reg}==18'b010101100000010111)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010101100000011000)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010101100000011001)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010101100000011010)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b010101100000011011)) color_data = 12'b011111001111;
		if(({row_reg, col_reg}>=18'b010101100000011100) && ({row_reg, col_reg}<18'b010101100000011110)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}>=18'b010101100000011110) && ({row_reg, col_reg}<18'b010101100000100000)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b010101100000100000)) color_data = 12'b010010011100;
		if(({row_reg, col_reg}==18'b010101100000100001)) color_data = 12'b001001111010;
		if(({row_reg, col_reg}>=18'b010101100000100010) && ({row_reg, col_reg}<18'b010101100000100100)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b010101100000100100)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010101100000100101)) color_data = 12'b000101111100;
		if(({row_reg, col_reg}>=18'b010101100000100110) && ({row_reg, col_reg}<18'b010101100000101010)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010101100000101010)) color_data = 12'b000101111100;
		if(({row_reg, col_reg}==18'b010101100000101011)) color_data = 12'b000101111011;
		if(({row_reg, col_reg}==18'b010101100000101100)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b010101100000101101)) color_data = 12'b001101111010;
		if(({row_reg, col_reg}==18'b010101100000101110)) color_data = 12'b001101111001;
		if(({row_reg, col_reg}==18'b010101100000101111)) color_data = 12'b010001101001;
		if(({row_reg, col_reg}>=18'b010101100000110000) && ({row_reg, col_reg}<18'b010101100000110010)) color_data = 12'b010101100111;
		if(({row_reg, col_reg}==18'b010101100000110010)) color_data = 12'b010101100110;
		if(({row_reg, col_reg}==18'b010101100000110011)) color_data = 12'b010101100111;
		if(({row_reg, col_reg}==18'b010101100000110100)) color_data = 12'b010001100110;
		if(({row_reg, col_reg}==18'b010101100000110101)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}>=18'b010101100000110110) && ({row_reg, col_reg}<18'b010101100000111010)) color_data = 12'b010101110111;
		if(({row_reg, col_reg}==18'b010101100000111010)) color_data = 12'b010101100110;
		if(({row_reg, col_reg}==18'b010101100000111011)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}==18'b010101100000111100)) color_data = 12'b010101100111;
		if(({row_reg, col_reg}==18'b010101100000111101)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}>=18'b010101100000111110) && ({row_reg, col_reg}<18'b010101100001000000)) color_data = 12'b010101100111;
		if(({row_reg, col_reg}==18'b010101100001000000)) color_data = 12'b010101110111;
		if(({row_reg, col_reg}==18'b010101100001000001)) color_data = 12'b010101100111;
		if(({row_reg, col_reg}==18'b010101100001000010)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==18'b010101100001000011)) color_data = 12'b010101100111;
		if(({row_reg, col_reg}==18'b010101100001000100)) color_data = 12'b010101100110;
		if(({row_reg, col_reg}>=18'b010101100001000101) && ({row_reg, col_reg}<18'b010101100001001010)) color_data = 12'b010101110111;
		if(({row_reg, col_reg}==18'b010101100001001010)) color_data = 12'b010001110111;
		if(({row_reg, col_reg}==18'b010101100001001011)) color_data = 12'b100111011110;
		if(({row_reg, col_reg}==18'b010101100001001100)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010101100001001101)) color_data = 12'b100011111110;
		if(({row_reg, col_reg}==18'b010101100001001110)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010101100001001111)) color_data = 12'b011011011110;
		if(({row_reg, col_reg}>=18'b010101100001010000) && ({row_reg, col_reg}<18'b010101100001010010)) color_data = 12'b000110001010;
		if(({row_reg, col_reg}==18'b010101100001010010)) color_data = 12'b000101111011;
		if(({row_reg, col_reg}==18'b010101100001010011)) color_data = 12'b000101111100;
		if(({row_reg, col_reg}==18'b010101100001010100)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b010101100001010101)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010101100001010110)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010101100001010111)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b010101100001011000)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}==18'b010101100001011001)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b010101100001011010)) color_data = 12'b000101111011;
		if(({row_reg, col_reg}>=18'b010101100001011011) && ({row_reg, col_reg}<18'b010101100001011101)) color_data = 12'b001001111010;
		if(({row_reg, col_reg}==18'b010101100001011101)) color_data = 12'b010010001011;
		if(({row_reg, col_reg}==18'b010101100001011110)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b010101100001011111)) color_data = 12'b101010111100;
		if(({row_reg, col_reg}==18'b010101100001100000)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}>=18'b010101100001100001) && ({row_reg, col_reg}<18'b010101100001100100)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010101100001100100)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==18'b010101100001100101)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010101100001100110)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==18'b010101100001100111)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010101100001101000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010101100001101001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010101100001101010)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010101100001101011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010101100001101100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010101100001101101) && ({row_reg, col_reg}<18'b010101100001110000)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==18'b010101100001110000)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010101100001110001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b010101100001110010) && ({row_reg, col_reg}<18'b010101100001110101)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010101100001110101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010101100001110110)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==18'b010101100001110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010101100001111000)) color_data = 12'b101010111010;
		if(({row_reg, col_reg}==18'b010101100001111001)) color_data = 12'b100110111010;
		if(({row_reg, col_reg}==18'b010101100001111010)) color_data = 12'b101011001011;
		if(({row_reg, col_reg}==18'b010101100001111011)) color_data = 12'b110011111101;
		if(({row_reg, col_reg}==18'b010101100001111100)) color_data = 12'b101111111101;
		if(({row_reg, col_reg}==18'b010101100001111101)) color_data = 12'b101011111110;
		if(({row_reg, col_reg}==18'b010101100001111110)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}==18'b010101100001111111)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010101100010000000) && ({row_reg, col_reg}<18'b010101100010000100)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010101100010000100)) color_data = 12'b010010101101;
		if(({row_reg, col_reg}==18'b010101100010000101)) color_data = 12'b000101101011;
		if(({row_reg, col_reg}==18'b010101100010000110)) color_data = 12'b001001101100;
		if(({row_reg, col_reg}==18'b010101100010000111)) color_data = 12'b001101101011;
		if(({row_reg, col_reg}==18'b010101100010001000)) color_data = 12'b010101111011;
		if(({row_reg, col_reg}==18'b010101100010001001)) color_data = 12'b010001101000;
		if(({row_reg, col_reg}==18'b010101100010001010)) color_data = 12'b010101111000;
		if(({row_reg, col_reg}>=18'b010101100010001011) && ({row_reg, col_reg}<18'b010101100010001110)) color_data = 12'b010101100111;
		if(({row_reg, col_reg}==18'b010101100010001110)) color_data = 12'b010101110111;
		if(({row_reg, col_reg}>=18'b010101100010001111) && ({row_reg, col_reg}<18'b010101100010010001)) color_data = 12'b010101100110;
		if(({row_reg, col_reg}==18'b010101100010010001)) color_data = 12'b010101110111;
		if(({row_reg, col_reg}>=18'b010101100010010010) && ({row_reg, col_reg}<18'b010101100010010100)) color_data = 12'b010101100111;
		if(({row_reg, col_reg}==18'b010101100010010100)) color_data = 12'b011001111000;
		if(({row_reg, col_reg}>=18'b010101100010010101) && ({row_reg, col_reg}<18'b010101100010011000)) color_data = 12'b011001101000;
		if(({row_reg, col_reg}>=18'b010101100010011000) && ({row_reg, col_reg}<18'b010101100010011010)) color_data = 12'b011001111000;
		if(({row_reg, col_reg}==18'b010101100010011010)) color_data = 12'b011001101000;
		if(({row_reg, col_reg}==18'b010101100010011011)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==18'b010101100010011100)) color_data = 12'b011001111000;
		if(({row_reg, col_reg}==18'b010101100010011101)) color_data = 12'b010101110111;
		if(({row_reg, col_reg}==18'b010101100010011110)) color_data = 12'b010101100111;
		if(({row_reg, col_reg}==18'b010101100010011111)) color_data = 12'b010001100110;
		if(({row_reg, col_reg}==18'b010101100010100000)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==18'b010101100010100001)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==18'b010101100010100010)) color_data = 12'b100110111011;
		if(({row_reg, col_reg}>=18'b010101100010100011) && ({row_reg, col_reg}<18'b010101100010100110)) color_data = 12'b100110101010;
		if(({row_reg, col_reg}==18'b010101100010100110)) color_data = 12'b100110111011;
		if(({row_reg, col_reg}>=18'b010101100010100111) && ({row_reg, col_reg}<18'b010101100010101001)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b010101100010101001)) color_data = 12'b101010111100;
		if(({row_reg, col_reg}==18'b010101100010101010)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}>=18'b010101100010101011) && ({row_reg, col_reg}<18'b010101100010101101)) color_data = 12'b101010101100;
		if(({row_reg, col_reg}==18'b010101100010101101)) color_data = 12'b100110111101;
		if(({row_reg, col_reg}==18'b010101100010101110)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b010101100010101111)) color_data = 12'b010110001011;
		if(({row_reg, col_reg}>=18'b010101100010110000) && ({row_reg, col_reg}<18'b010101100010110010)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010101100010110010)) color_data = 12'b001101111011;
		if(({row_reg, col_reg}==18'b010101100010110011)) color_data = 12'b010001111010;
		if(({row_reg, col_reg}==18'b010101100010110100)) color_data = 12'b010101111001;
		if(({row_reg, col_reg}==18'b010101100010110101)) color_data = 12'b010101111000;
		if(({row_reg, col_reg}==18'b010101100010110110)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}>=18'b010101100010110111) && ({row_reg, col_reg}<18'b010101100010111010)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}==18'b010101100010111010)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}==18'b010101100010111011)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010101100010111100) && ({row_reg, col_reg}<18'b010101100011000000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010101100011000000) && ({row_reg, col_reg}<18'b010101100011001111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010101100011001111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010101100011010000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010101100011010001) && ({row_reg, col_reg}<18'b010101100011010101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010101100011010101)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010101100011010110) && ({row_reg, col_reg}<18'b010101100011110101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010101100011110101)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}==18'b010101100011110110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010101100011110111)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}==18'b010101100011111000)) color_data = 12'b010101100110;
		if(({row_reg, col_reg}==18'b010101100011111001)) color_data = 12'b010101110111;
		if(({row_reg, col_reg}==18'b010101100011111010)) color_data = 12'b010001111000;
		if(({row_reg, col_reg}==18'b010101100011111011)) color_data = 12'b100011001101;
		if(({row_reg, col_reg}==18'b010101100011111100)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}>=18'b010101100011111101) && ({row_reg, col_reg}<18'b010101100011111111)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010101100011111111) && ({row_reg, col_reg}<18'b010101100100000001)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010101100100000001)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010101100100000010)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010101100100000011)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010101100100000100)) color_data = 12'b011111011110;
		if(({row_reg, col_reg}==18'b010101100100000101)) color_data = 12'b011011001101;
		if(({row_reg, col_reg}==18'b010101100100000110)) color_data = 12'b010110111100;
		if(({row_reg, col_reg}>=18'b010101100100000111) && ({row_reg, col_reg}<18'b010101100100001001)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}==18'b010101100100001001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010101100100001010)) color_data = 12'b011010101101;

		if(({row_reg, col_reg}>=18'b010101100100001011) && ({row_reg, col_reg}<18'b010101101000000000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010101101000000000)) color_data = 12'b010010011101;
		if(({row_reg, col_reg}==18'b010101101000000001)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}==18'b010101101000000010)) color_data = 12'b010010001110;
		if(({row_reg, col_reg}==18'b010101101000000011)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}>=18'b010101101000000100) && ({row_reg, col_reg}<18'b010101101000000110)) color_data = 12'b010010001110;
		if(({row_reg, col_reg}==18'b010101101000000110)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}==18'b010101101000000111)) color_data = 12'b010110001101;
		if(({row_reg, col_reg}>=18'b010101101000001000) && ({row_reg, col_reg}<18'b010101101000001110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010101101000001110) && ({row_reg, col_reg}<18'b010101101000010000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010101101000010000) && ({row_reg, col_reg}<18'b010101101000010100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010101101000010100)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b010101101000010101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010101101000010110)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}>=18'b010101101000010111) && ({row_reg, col_reg}<18'b010101101000011001)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}==18'b010101101000011001)) color_data = 12'b010010011101;
		if(({row_reg, col_reg}==18'b010101101000011010)) color_data = 12'b010010001100;
		if(({row_reg, col_reg}==18'b010101101000011011)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==18'b010101101000011100)) color_data = 12'b100011001111;
		if(({row_reg, col_reg}==18'b010101101000011101)) color_data = 12'b100011011111;
		if(({row_reg, col_reg}==18'b010101101000011110)) color_data = 12'b011111001111;
		if(({row_reg, col_reg}==18'b010101101000011111)) color_data = 12'b100011011111;
		if(({row_reg, col_reg}==18'b010101101000100000)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}>=18'b010101101000100001) && ({row_reg, col_reg}<18'b010101101000100100)) color_data = 12'b010110111101;
		if(({row_reg, col_reg}>=18'b010101101000100100) && ({row_reg, col_reg}<18'b010101101000101100)) color_data = 12'b010110111110;
		if(({row_reg, col_reg}==18'b010101101000101100)) color_data = 12'b010110111101;
		if(({row_reg, col_reg}==18'b010101101000101101)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}==18'b010101101000101110)) color_data = 12'b011010101100;
		if(({row_reg, col_reg}==18'b010101101000101111)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}>=18'b010101101000110000) && ({row_reg, col_reg}<18'b010101101000110010)) color_data = 12'b011110101011;
		if(({row_reg, col_reg}==18'b010101101000110010)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}==18'b010101101000110011)) color_data = 12'b011110011001;
		if(({row_reg, col_reg}==18'b010101101000110100)) color_data = 12'b011010001001;
		if(({row_reg, col_reg}==18'b010101101000110101)) color_data = 12'b011010011010;
		if(({row_reg, col_reg}==18'b010101101000110110)) color_data = 12'b011010001001;
		if(({row_reg, col_reg}==18'b010101101000110111)) color_data = 12'b010110001001;
		if(({row_reg, col_reg}==18'b010101101000111000)) color_data = 12'b011110011010;
		if(({row_reg, col_reg}==18'b010101101000111001)) color_data = 12'b011110101010;
		if(({row_reg, col_reg}>=18'b010101101000111010) && ({row_reg, col_reg}<18'b010101101000111100)) color_data = 12'b011110011010;
		if(({row_reg, col_reg}==18'b010101101000111100)) color_data = 12'b011110101011;
		if(({row_reg, col_reg}==18'b010101101000111101)) color_data = 12'b011110011010;
		if(({row_reg, col_reg}>=18'b010101101000111110) && ({row_reg, col_reg}<18'b010101101001000000)) color_data = 12'b011010001001;
		if(({row_reg, col_reg}==18'b010101101001000000)) color_data = 12'b011010011001;
		if(({row_reg, col_reg}==18'b010101101001000001)) color_data = 12'b011110011010;
		if(({row_reg, col_reg}>=18'b010101101001000010) && ({row_reg, col_reg}<18'b010101101001000101)) color_data = 12'b011110101010;
		if(({row_reg, col_reg}==18'b010101101001000101)) color_data = 12'b011110101011;
		if(({row_reg, col_reg}>=18'b010101101001000110) && ({row_reg, col_reg}<18'b010101101001001001)) color_data = 12'b011110101010;
		if(({row_reg, col_reg}>=18'b010101101001001001) && ({row_reg, col_reg}<18'b010101101001001011)) color_data = 12'b011010101010;
		if(({row_reg, col_reg}==18'b010101101001001011)) color_data = 12'b100011101110;
		if(({row_reg, col_reg}==18'b010101101001001100)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010101101001001101) && ({row_reg, col_reg}<18'b010101101001001111)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010101101001001111)) color_data = 12'b011111101111;
		if(({row_reg, col_reg}>=18'b010101101001010000) && ({row_reg, col_reg}<18'b010101101001010010)) color_data = 12'b010110111101;
		if(({row_reg, col_reg}==18'b010101101001010010)) color_data = 12'b010010111101;
		if(({row_reg, col_reg}==18'b010101101001010011)) color_data = 12'b010010111110;
		if(({row_reg, col_reg}==18'b010101101001010100)) color_data = 12'b010010011110;
		if(({row_reg, col_reg}==18'b010101101001010101)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010101101001010110)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b010101101001010111)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}==18'b010101101001011000)) color_data = 12'b001010001110;
		if(({row_reg, col_reg}==18'b010101101001011001)) color_data = 12'b010010011110;
		if(({row_reg, col_reg}>=18'b010101101001011010) && ({row_reg, col_reg}<18'b010101101001011100)) color_data = 12'b010110111101;
		if(({row_reg, col_reg}==18'b010101101001011100)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}==18'b010101101001011101)) color_data = 12'b011110111101;
		if(({row_reg, col_reg}==18'b010101101001011110)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b010101101001011111)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}>=18'b010101101001100000) && ({row_reg, col_reg}<18'b010101101001100011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010101101001100011)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b010101101001100100) && ({row_reg, col_reg}<18'b010101101001100110)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==18'b010101101001100110)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010101101001100111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b010101101001101000) && ({row_reg, col_reg}<18'b010101101001101100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}>=18'b010101101001101100) && ({row_reg, col_reg}<18'b010101101001101110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010101101001101110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010101101001101111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010101101001110000)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==18'b010101101001110001)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==18'b010101101001110010)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}>=18'b010101101001110011) && ({row_reg, col_reg}<18'b010101101001110110)) color_data = 12'b100110001000;
		if(({row_reg, col_reg}==18'b010101101001110110)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010101101001110111)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010101101001111000)) color_data = 12'b101010111010;
		if(({row_reg, col_reg}==18'b010101101001111001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010101101001111010)) color_data = 12'b101010111010;
		if(({row_reg, col_reg}==18'b010101101001111011)) color_data = 12'b101011001011;
		if(({row_reg, col_reg}==18'b010101101001111100)) color_data = 12'b100111001011;
		if(({row_reg, col_reg}==18'b010101101001111101)) color_data = 12'b100111011101;
		if(({row_reg, col_reg}==18'b010101101001111110)) color_data = 12'b100011011110;
		if(({row_reg, col_reg}==18'b010101101001111111)) color_data = 12'b011111001110;
		if(({row_reg, col_reg}>=18'b010101101010000000) && ({row_reg, col_reg}<18'b010101101010000011)) color_data = 12'b011011001110;
		if(({row_reg, col_reg}>=18'b010101101010000011) && ({row_reg, col_reg}<18'b010101101010000101)) color_data = 12'b010111001110;
		if(({row_reg, col_reg}==18'b010101101010000101)) color_data = 12'b010110111110;
		if(({row_reg, col_reg}==18'b010101101010000110)) color_data = 12'b011010111111;
		if(({row_reg, col_reg}==18'b010101101010000111)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==18'b010101101010001000)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}>=18'b010101101010001001) && ({row_reg, col_reg}<18'b010101101010001011)) color_data = 12'b010001111010;
		if(({row_reg, col_reg}==18'b010101101010001011)) color_data = 12'b010110001010;
		if(({row_reg, col_reg}==18'b010101101010001100)) color_data = 12'b010001111001;
		if(({row_reg, col_reg}==18'b010101101010001101)) color_data = 12'b010110001010;
		if(({row_reg, col_reg}>=18'b010101101010001110) && ({row_reg, col_reg}<18'b010101101010010001)) color_data = 12'b011110101010;
		if(({row_reg, col_reg}==18'b010101101010010001)) color_data = 12'b011110101011;
		if(({row_reg, col_reg}==18'b010101101010010010)) color_data = 12'b011010011010;
		if(({row_reg, col_reg}==18'b010101101010010011)) color_data = 12'b010001111001;
		if(({row_reg, col_reg}>=18'b010101101010010100) && ({row_reg, col_reg}<18'b010101101010011010)) color_data = 12'b010101111010;
		if(({row_reg, col_reg}==18'b010101101010011010)) color_data = 12'b010001111001;
		if(({row_reg, col_reg}==18'b010101101010011011)) color_data = 12'b010001111000;
		if(({row_reg, col_reg}==18'b010101101010011100)) color_data = 12'b011110101011;
		if(({row_reg, col_reg}==18'b010101101010011101)) color_data = 12'b011110101010;
		if(({row_reg, col_reg}>=18'b010101101010011110) && ({row_reg, col_reg}<18'b010101101010100000)) color_data = 12'b011010101010;
		if(({row_reg, col_reg}==18'b010101101010100000)) color_data = 12'b100010101010;
		if(({row_reg, col_reg}>=18'b010101101010100001) && ({row_reg, col_reg}<18'b010101101010100111)) color_data = 12'b100111001100;
		if(({row_reg, col_reg}==18'b010101101010100111)) color_data = 12'b100011001100;
		if(({row_reg, col_reg}==18'b010101101010101000)) color_data = 12'b100111001100;
		if(({row_reg, col_reg}==18'b010101101010101001)) color_data = 12'b100111001101;
		if(({row_reg, col_reg}==18'b010101101010101010)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}==18'b010101101010101011)) color_data = 12'b011110011011;
		if(({row_reg, col_reg}==18'b010101101010101100)) color_data = 12'b011110011100;
		if(({row_reg, col_reg}==18'b010101101010101101)) color_data = 12'b011110011101;
		if(({row_reg, col_reg}==18'b010101101010101110)) color_data = 12'b011010011100;
		if(({row_reg, col_reg}==18'b010101101010101111)) color_data = 12'b010010001011;
		if(({row_reg, col_reg}==18'b010101101010110000)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010101101010110001)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b010101101010110010)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}>=18'b010101101010110011) && ({row_reg, col_reg}<18'b010101101010110101)) color_data = 12'b010001111011;
		if(({row_reg, col_reg}==18'b010101101010110101)) color_data = 12'b010001111010;
		if(({row_reg, col_reg}==18'b010101101010110110)) color_data = 12'b010101111001;
		if(({row_reg, col_reg}==18'b010101101010110111)) color_data = 12'b011001111001;
		if(({row_reg, col_reg}==18'b010101101010111000)) color_data = 12'b011001111000;
		if(({row_reg, col_reg}==18'b010101101010111001)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==18'b010101101010111010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010101101010111011) && ({row_reg, col_reg}<18'b010101101010111101)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}==18'b010101101010111101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010101101010111110) && ({row_reg, col_reg}<18'b010101101011000000)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010101101011000000) && ({row_reg, col_reg}<18'b010101101011010000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010101101011010000)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010101101011010001) && ({row_reg, col_reg}<18'b010101101011010100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010101101011010100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010101101011010101) && ({row_reg, col_reg}<18'b010101101011110011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010101101011110011)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==18'b010101101011110100)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==18'b010101101011110101)) color_data = 12'b010101100110;
		if(({row_reg, col_reg}==18'b010101101011110110)) color_data = 12'b011110001000;
		if(({row_reg, col_reg}==18'b010101101011110111)) color_data = 12'b100010101010;
		if(({row_reg, col_reg}==18'b010101101011111000)) color_data = 12'b011110011001;
		if(({row_reg, col_reg}==18'b010101101011111001)) color_data = 12'b011110011010;
		if(({row_reg, col_reg}==18'b010101101011111010)) color_data = 12'b011010011010;
		if(({row_reg, col_reg}==18'b010101101011111011)) color_data = 12'b011110111101;
		if(({row_reg, col_reg}>=18'b010101101011111100) && ({row_reg, col_reg}<18'b010101101011111111)) color_data = 12'b011011001110;
		if(({row_reg, col_reg}==18'b010101101011111111)) color_data = 12'b010111001110;
		if(({row_reg, col_reg}>=18'b010101101100000000) && ({row_reg, col_reg}<18'b010101101100000011)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010101101100000011)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010101101100000100)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010101101100000101)) color_data = 12'b011111011110;
		if(({row_reg, col_reg}==18'b010101101100000110)) color_data = 12'b011011011110;
		if(({row_reg, col_reg}>=18'b010101101100000111) && ({row_reg, col_reg}<18'b010101101100001001)) color_data = 12'b011111011110;
		if(({row_reg, col_reg}==18'b010101101100001001)) color_data = 12'b011111001110;
		if(({row_reg, col_reg}==18'b010101101100001010)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==18'b010101101100001011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010101101100001100)) color_data = 12'b011010101111;

		if(({row_reg, col_reg}>=18'b010101101100001101) && ({row_reg, col_reg}<18'b010101110000000000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010101110000000000)) color_data = 12'b011010111111;
		if(({row_reg, col_reg}>=18'b010101110000000001) && ({row_reg, col_reg}<18'b010101110000001001)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b010101110000001001)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}>=18'b010101110000001010) && ({row_reg, col_reg}<18'b010101110000001100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010101110000001100) && ({row_reg, col_reg}<18'b010101110000001110)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b010101110000001110)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}==18'b010101110000001111)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b010101110000010000) && ({row_reg, col_reg}<18'b010101110000011000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010101110000011000)) color_data = 12'b011010111111;
		if(({row_reg, col_reg}==18'b010101110000011001)) color_data = 12'b011110111111;
		if(({row_reg, col_reg}==18'b010101110000011010)) color_data = 12'b011010111111;
		if(({row_reg, col_reg}>=18'b010101110000011011) && ({row_reg, col_reg}<18'b010101110000011101)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==18'b010101110000011101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010101110000011110)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}==18'b010101110000011111)) color_data = 12'b011110111110;
		if(({row_reg, col_reg}==18'b010101110000100000)) color_data = 12'b100011011111;
		if(({row_reg, col_reg}>=18'b010101110000100001) && ({row_reg, col_reg}<18'b010101110000100011)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}>=18'b010101110000100011) && ({row_reg, col_reg}<18'b010101110000101110)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010101110000101110)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}==18'b010101110000101111)) color_data = 12'b101011101111;
		if(({row_reg, col_reg}>=18'b010101110000110000) && ({row_reg, col_reg}<18'b010101110000110011)) color_data = 12'b101111101111;
		if(({row_reg, col_reg}==18'b010101110000110011)) color_data = 12'b100010111101;
		if(({row_reg, col_reg}>=18'b010101110000110100) && ({row_reg, col_reg}<18'b010101110000110111)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}==18'b010101110000110111)) color_data = 12'b100010111101;
		if(({row_reg, col_reg}==18'b010101110000111000)) color_data = 12'b101011101111;
		if(({row_reg, col_reg}==18'b010101110000111001)) color_data = 12'b101111101111;
		if(({row_reg, col_reg}==18'b010101110000111010)) color_data = 12'b101111111111;
		if(({row_reg, col_reg}==18'b010101110000111011)) color_data = 12'b101111101111;
		if(({row_reg, col_reg}==18'b010101110000111100)) color_data = 12'b101011011111;
		if(({row_reg, col_reg}==18'b010101110000111101)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}>=18'b010101110000111110) && ({row_reg, col_reg}<18'b010101110001000001)) color_data = 12'b011010101011;
		if(({row_reg, col_reg}==18'b010101110001000001)) color_data = 12'b100111011110;
		if(({row_reg, col_reg}==18'b010101110001000010)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}>=18'b010101110001000011) && ({row_reg, col_reg}<18'b010101110001000101)) color_data = 12'b101011111110;
		if(({row_reg, col_reg}>=18'b010101110001000101) && ({row_reg, col_reg}<18'b010101110001001000)) color_data = 12'b101011101111;
		if(({row_reg, col_reg}>=18'b010101110001001000) && ({row_reg, col_reg}<18'b010101110001001010)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}==18'b010101110001001010)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010101110001001011) && ({row_reg, col_reg}<18'b010101110001001101)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010101110001001101)) color_data = 12'b011111111111;
		if(({row_reg, col_reg}>=18'b010101110001001110) && ({row_reg, col_reg}<18'b010101110001010000)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010101110001010000)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}>=18'b010101110001010001) && ({row_reg, col_reg}<18'b010101110001010011)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010101110001010011)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010101110001010100)) color_data = 12'b011011001111;
		if(({row_reg, col_reg}==18'b010101110001010101)) color_data = 12'b000101111011;
		if(({row_reg, col_reg}==18'b010101110001010110)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010101110001010111)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b010101110001011000)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010101110001011001)) color_data = 12'b011011001111;
		if(({row_reg, col_reg}>=18'b010101110001011010) && ({row_reg, col_reg}<18'b010101110001011100)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010101110001011100)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}==18'b010101110001011101)) color_data = 12'b101011011111;
		if(({row_reg, col_reg}==18'b010101110001011110)) color_data = 12'b100110111100;
		if(({row_reg, col_reg}==18'b010101110001011111)) color_data = 12'b100110111011;
		if(({row_reg, col_reg}>=18'b010101110001100000) && ({row_reg, col_reg}<18'b010101110001100011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010101110001100011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010101110001100100) && ({row_reg, col_reg}<18'b010101110001100111)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b010101110001100111) && ({row_reg, col_reg}<18'b010101110001101010)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010101110001101010) && ({row_reg, col_reg}<18'b010101110001101100)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==18'b010101110001101100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010101110001101101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010101110001101110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010101110001101111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010101110001110000)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==18'b010101110001110001)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010101110001110010)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b010101110001110011) && ({row_reg, col_reg}<18'b010101110001110101)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==18'b010101110001110101)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==18'b010101110001110110)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==18'b010101110001110111)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010101110001111000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}==18'b010101110001111001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010101110001111010) && ({row_reg, col_reg}<18'b010101110001111100)) color_data = 12'b101010111011;
		if(({row_reg, col_reg}==18'b010101110001111100)) color_data = 12'b100110111010;
		if(({row_reg, col_reg}==18'b010101110001111101)) color_data = 12'b100010111100;
		if(({row_reg, col_reg}==18'b010101110001111110)) color_data = 12'b011110111100;
		if(({row_reg, col_reg}==18'b010101110001111111)) color_data = 12'b010110011011;
		if(({row_reg, col_reg}>=18'b010101110010000000) && ({row_reg, col_reg}<18'b010101110010000010)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}>=18'b010101110010000010) && ({row_reg, col_reg}<18'b010101110010000100)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b010101110010000100)) color_data = 12'b011011011111;
		if(({row_reg, col_reg}==18'b010101110010000101)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010101110010000110) && ({row_reg, col_reg}<18'b010101110010001000)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010101110010001000)) color_data = 12'b100011011111;
		if(({row_reg, col_reg}==18'b010101110010001001)) color_data = 12'b010010001100;
		if(({row_reg, col_reg}>=18'b010101110010001010) && ({row_reg, col_reg}<18'b010101110010001100)) color_data = 12'b001101111011;
		if(({row_reg, col_reg}==18'b010101110010001100)) color_data = 12'b001101111010;
		if(({row_reg, col_reg}==18'b010101110010001101)) color_data = 12'b011010101100;
		if(({row_reg, col_reg}==18'b010101110010001110)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}==18'b010101110010001111)) color_data = 12'b101111111111;
		if(({row_reg, col_reg}>=18'b010101110010010000) && ({row_reg, col_reg}<18'b010101110010010010)) color_data = 12'b101011101111;
		if(({row_reg, col_reg}==18'b010101110010010010)) color_data = 12'b011110111101;
		if(({row_reg, col_reg}==18'b010101110010010011)) color_data = 12'b001101111010;
		if(({row_reg, col_reg}==18'b010101110010010100)) color_data = 12'b001101111011;
		if(({row_reg, col_reg}>=18'b010101110010010101) && ({row_reg, col_reg}<18'b010101110010011000)) color_data = 12'b010001111100;
		if(({row_reg, col_reg}>=18'b010101110010011000) && ({row_reg, col_reg}<18'b010101110010011010)) color_data = 12'b010001111011;
		if(({row_reg, col_reg}==18'b010101110010011010)) color_data = 12'b010001111010;
		if(({row_reg, col_reg}==18'b010101110010011011)) color_data = 12'b010010011010;
		if(({row_reg, col_reg}==18'b010101110010011100)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}>=18'b010101110010011101) && ({row_reg, col_reg}<18'b010101110010100010)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}>=18'b010101110010100010) && ({row_reg, col_reg}<18'b010101110010100100)) color_data = 12'b101011111110;
		if(({row_reg, col_reg}==18'b010101110010100100)) color_data = 12'b100111101110;
		if(({row_reg, col_reg}>=18'b010101110010100101) && ({row_reg, col_reg}<18'b010101110010100111)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}>=18'b010101110010100111) && ({row_reg, col_reg}<18'b010101110010101010)) color_data = 12'b100111101110;
		if(({row_reg, col_reg}==18'b010101110010101010)) color_data = 12'b011010101011;
		if(({row_reg, col_reg}==18'b010101110010101011)) color_data = 12'b001101111010;
		if(({row_reg, col_reg}==18'b010101110010101100)) color_data = 12'b001101111011;
		if(({row_reg, col_reg}==18'b010101110010101101)) color_data = 12'b010001111011;
		if(({row_reg, col_reg}==18'b010101110010101110)) color_data = 12'b001101111011;
		if(({row_reg, col_reg}==18'b010101110010101111)) color_data = 12'b001001111010;
		if(({row_reg, col_reg}>=18'b010101110010110000) && ({row_reg, col_reg}<18'b010101110010110010)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b010101110010110010) && ({row_reg, col_reg}<18'b010101110010110100)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}>=18'b010101110010110100) && ({row_reg, col_reg}<18'b010101110010110110)) color_data = 12'b010001111100;
		if(({row_reg, col_reg}==18'b010101110010110110)) color_data = 12'b010101111100;
		if(({row_reg, col_reg}==18'b010101110010110111)) color_data = 12'b010101111011;
		if(({row_reg, col_reg}==18'b010101110010111000)) color_data = 12'b011001111001;
		if(({row_reg, col_reg}==18'b010101110010111001)) color_data = 12'b011001111000;
		if(({row_reg, col_reg}==18'b010101110010111010)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}>=18'b010101110010111011) && ({row_reg, col_reg}<18'b010101110010111110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010101110010111110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010101110010111111) && ({row_reg, col_reg}<18'b010101110011000001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010101110011000001) && ({row_reg, col_reg}<18'b010101110011010001)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010101110011010001) && ({row_reg, col_reg}<18'b010101110011010011)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010101110011010011) && ({row_reg, col_reg}<18'b010101110011101100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010101110011101100)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010101110011101101) && ({row_reg, col_reg}<18'b010101110011101111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010101110011101111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010101110011110000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010101110011110001) && ({row_reg, col_reg}<18'b010101110011110011)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010101110011110011) && ({row_reg, col_reg}<18'b010101110011110101)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==18'b010101110011110101)) color_data = 12'b010101100111;
		if(({row_reg, col_reg}==18'b010101110011110110)) color_data = 12'b100010101010;
		if(({row_reg, col_reg}==18'b010101110011110111)) color_data = 12'b110011101110;
		if(({row_reg, col_reg}==18'b010101110011111000)) color_data = 12'b110011111110;
		if(({row_reg, col_reg}==18'b010101110011111001)) color_data = 12'b101111101110;
		if(({row_reg, col_reg}==18'b010101110011111010)) color_data = 12'b101111111111;
		if(({row_reg, col_reg}==18'b010101110011111011)) color_data = 12'b010110101100;
		if(({row_reg, col_reg}==18'b010101110011111100)) color_data = 12'b001001111010;
		if(({row_reg, col_reg}==18'b010101110011111101)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}>=18'b010101110011111110) && ({row_reg, col_reg}<18'b010101110100000000)) color_data = 12'b000110001011;
		if(({row_reg, col_reg}==18'b010101110100000000)) color_data = 12'b011111101110;
		if(({row_reg, col_reg}==18'b010101110100000001)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010101110100000010) && ({row_reg, col_reg}<18'b010101110100000101)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010101110100000101) && ({row_reg, col_reg}<18'b010101110100000111)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010101110100000111) && ({row_reg, col_reg}<18'b010101110100001001)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010101110100001001)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}==18'b010101110100001010)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==18'b010101110100001011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010101110100001100)) color_data = 12'b011010101111;

		if(({row_reg, col_reg}>=18'b010101110100001101) && ({row_reg, col_reg}<18'b010101111000000000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010101111000000000)) color_data = 12'b011110111111;
		if(({row_reg, col_reg}>=18'b010101111000000001) && ({row_reg, col_reg}<18'b010101111000001000)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b010101111000001000) && ({row_reg, col_reg}<18'b010101111000001010)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}>=18'b010101111000001010) && ({row_reg, col_reg}<18'b010101111000010000)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b010101111000010000) && ({row_reg, col_reg}<18'b010101111000011111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010101111000011111)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==18'b010101111000100000)) color_data = 12'b100011011111;
		if(({row_reg, col_reg}==18'b010101111000100001)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010101111000100010)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b010101111000100011)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010101111000100100) && ({row_reg, col_reg}<18'b010101111000101001)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010101111000101001) && ({row_reg, col_reg}<18'b010101111000101111)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010101111000101111)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}>=18'b010101111000110000) && ({row_reg, col_reg}<18'b010101111000110011)) color_data = 12'b101011101111;
		if(({row_reg, col_reg}==18'b010101111000110011)) color_data = 12'b100010111101;
		if(({row_reg, col_reg}==18'b010101111000110100)) color_data = 12'b011110101100;
		if(({row_reg, col_reg}==18'b010101111000110101)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b010101111000110110)) color_data = 12'b011010101100;
		if(({row_reg, col_reg}==18'b010101111000110111)) color_data = 12'b100010111101;
		if(({row_reg, col_reg}>=18'b010101111000111000) && ({row_reg, col_reg}<18'b010101111000111100)) color_data = 12'b101011101111;
		if(({row_reg, col_reg}==18'b010101111000111100)) color_data = 12'b100111011110;
		if(({row_reg, col_reg}==18'b010101111000111101)) color_data = 12'b011010111100;
		if(({row_reg, col_reg}==18'b010101111000111110)) color_data = 12'b011110111101;
		if(({row_reg, col_reg}==18'b010101111000111111)) color_data = 12'b011110111100;
		if(({row_reg, col_reg}==18'b010101111001000000)) color_data = 12'b011010111011;
		if(({row_reg, col_reg}==18'b010101111001000001)) color_data = 12'b100011011110;
		if(({row_reg, col_reg}==18'b010101111001000010)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}>=18'b010101111001000011) && ({row_reg, col_reg}<18'b010101111001001010)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010101111001001010) && ({row_reg, col_reg}<18'b010101111001001100)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010101111001001100)) color_data = 12'b011111111111;
		if(({row_reg, col_reg}==18'b010101111001001101)) color_data = 12'b011111101110;
		if(({row_reg, col_reg}>=18'b010101111001001110) && ({row_reg, col_reg}<18'b010101111001010000)) color_data = 12'b011111111111;
		if(({row_reg, col_reg}>=18'b010101111001010000) && ({row_reg, col_reg}<18'b010101111001010100)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010101111001010100)) color_data = 12'b011011001111;
		if(({row_reg, col_reg}==18'b010101111001010101)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}>=18'b010101111001010110) && ({row_reg, col_reg}<18'b010101111001011000)) color_data = 12'b001010001101;
		if(({row_reg, col_reg}==18'b010101111001011000)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b010101111001011001)) color_data = 12'b011011011111;
		if(({row_reg, col_reg}==18'b010101111001011010)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010101111001011011)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010101111001011100)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b010101111001011101)) color_data = 12'b101011101111;
		if(({row_reg, col_reg}==18'b010101111001011110)) color_data = 12'b100111001100;
		if(({row_reg, col_reg}==18'b010101111001011111)) color_data = 12'b100110111010;
		if(({row_reg, col_reg}>=18'b010101111001100000) && ({row_reg, col_reg}<18'b010101111001100010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010101111001100010)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==18'b010101111001100011)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010101111001100100) && ({row_reg, col_reg}<18'b010101111001100111)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010101111001100111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010101111001101000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010101111001101001) && ({row_reg, col_reg}<18'b010101111001101011)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==18'b010101111001101011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010101111001101100)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}==18'b010101111001101101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010101111001101110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010101111001101111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010101111001110000)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}>=18'b010101111001110001) && ({row_reg, col_reg}<18'b010101111001110101)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==18'b010101111001110101)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}>=18'b010101111001110110) && ({row_reg, col_reg}<18'b010101111001111000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010101111001111000)) color_data = 12'b101110111011;
		if(({row_reg, col_reg}>=18'b010101111001111001) && ({row_reg, col_reg}<18'b010101111001111011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010101111001111011)) color_data = 12'b101010111011;
		if(({row_reg, col_reg}==18'b010101111001111100)) color_data = 12'b100110111011;
		if(({row_reg, col_reg}==18'b010101111001111101)) color_data = 12'b100110111100;
		if(({row_reg, col_reg}==18'b010101111001111110)) color_data = 12'b100010111101;
		if(({row_reg, col_reg}==18'b010101111001111111)) color_data = 12'b011010011100;
		if(({row_reg, col_reg}>=18'b010101111010000000) && ({row_reg, col_reg}<18'b010101111010000010)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010101111010000010)) color_data = 12'b001010001101;
		if(({row_reg, col_reg}==18'b010101111010000011)) color_data = 12'b001010011101;
		if(({row_reg, col_reg}==18'b010101111010000100)) color_data = 12'b011011011111;
		if(({row_reg, col_reg}==18'b010101111010000101)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010101111010000110)) color_data = 12'b100011111110;
		if(({row_reg, col_reg}==18'b010101111010000111)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010101111010001000)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010101111010001001)) color_data = 12'b010010011101;
		if(({row_reg, col_reg}==18'b010101111010001010)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010101111010001011)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b010101111010001100)) color_data = 12'b001001111010;
		if(({row_reg, col_reg}==18'b010101111010001101)) color_data = 12'b010110101100;
		if(({row_reg, col_reg}>=18'b010101111010001110) && ({row_reg, col_reg}<18'b010101111010010000)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b010101111010010000)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010101111010010001)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b010101111010010010)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}==18'b010101111010010011)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b010101111010010100)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}>=18'b010101111010010101) && ({row_reg, col_reg}<18'b010101111010011000)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010101111010011000)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010101111010011001)) color_data = 12'b001101111011;
		if(({row_reg, col_reg}==18'b010101111010011010)) color_data = 12'b001101111010;
		if(({row_reg, col_reg}==18'b010101111010011011)) color_data = 12'b001110011011;
		if(({row_reg, col_reg}==18'b010101111010011100)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010101111010011101)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010101111010011110)) color_data = 12'b100011101110;
		if(({row_reg, col_reg}>=18'b010101111010011111) && ({row_reg, col_reg}<18'b010101111010100010)) color_data = 12'b100111111110;
		if(({row_reg, col_reg}==18'b010101111010100010)) color_data = 12'b100011111110;
		if(({row_reg, col_reg}>=18'b010101111010100011) && ({row_reg, col_reg}<18'b010101111010100110)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010101111010100110)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}==18'b010101111010100111)) color_data = 12'b100111111110;
		if(({row_reg, col_reg}>=18'b010101111010101000) && ({row_reg, col_reg}<18'b010101111010101010)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010101111010101010)) color_data = 12'b010110101100;
		if(({row_reg, col_reg}==18'b010101111010101011)) color_data = 12'b001101111011;
		if(({row_reg, col_reg}>=18'b010101111010101100) && ({row_reg, col_reg}<18'b010101111010101110)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010101111010101110)) color_data = 12'b001101111011;
		if(({row_reg, col_reg}==18'b010101111010101111)) color_data = 12'b001110001011;
		if(({row_reg, col_reg}==18'b010101111010110000)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b010101111010110001)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010101111010110010) && ({row_reg, col_reg}<18'b010101111010110101)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010101111010110101)) color_data = 12'b010001111101;
		if(({row_reg, col_reg}==18'b010101111010110110)) color_data = 12'b010001101100;
		if(({row_reg, col_reg}==18'b010101111010110111)) color_data = 12'b010101111011;
		if(({row_reg, col_reg}==18'b010101111010111000)) color_data = 12'b010101111001;
		if(({row_reg, col_reg}==18'b010101111010111001)) color_data = 12'b010101110111;
		if(({row_reg, col_reg}>=18'b010101111010111010) && ({row_reg, col_reg}<18'b010101111010111100)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}==18'b010101111010111100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010101111010111101) && ({row_reg, col_reg}<18'b010101111011000000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010101111011000000) && ({row_reg, col_reg}<18'b010101111011110000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010101111011110000)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==18'b010101111011110001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010101111011110010) && ({row_reg, col_reg}<18'b010101111011110100)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}>=18'b010101111011110100) && ({row_reg, col_reg}<18'b010101111011110110)) color_data = 12'b010101110111;
		if(({row_reg, col_reg}==18'b010101111011110110)) color_data = 12'b100010101010;
		if(({row_reg, col_reg}>=18'b010101111011110111) && ({row_reg, col_reg}<18'b010101111011111001)) color_data = 12'b101111101110;
		if(({row_reg, col_reg}==18'b010101111011111001)) color_data = 12'b101011101110;
		if(({row_reg, col_reg}==18'b010101111011111010)) color_data = 12'b101011101111;
		if(({row_reg, col_reg}==18'b010101111011111011)) color_data = 12'b010110101100;
		if(({row_reg, col_reg}==18'b010101111011111100)) color_data = 12'b000101111010;
		if(({row_reg, col_reg}==18'b010101111011111101)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b010101111011111110)) color_data = 12'b000110001011;
		if(({row_reg, col_reg}==18'b010101111011111111)) color_data = 12'b000110011011;
		if(({row_reg, col_reg}==18'b010101111100000000)) color_data = 12'b100011101110;
		if(({row_reg, col_reg}==18'b010101111100000001)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010101111100000010)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010101111100000011)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010101111100000100) && ({row_reg, col_reg}<18'b010101111100001000)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010101111100001000)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010101111100001001)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}==18'b010101111100001010)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}>=18'b010101111100001011) && ({row_reg, col_reg}<18'b010101111100010000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010101111100010000)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b010101111100010001) && ({row_reg, col_reg}<18'b010110000000001111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010110000000001111)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010110000000010000) && ({row_reg, col_reg}<18'b010110000000010110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010110000000010110) && ({row_reg, col_reg}<18'b010110000000011110)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b010110000000011110) && ({row_reg, col_reg}<18'b010110000000100000)) color_data = 12'b011010111111;
		if(({row_reg, col_reg}==18'b010110000000100000)) color_data = 12'b100011101110;
		if(({row_reg, col_reg}>=18'b010110000000100001) && ({row_reg, col_reg}<18'b010110000000100101)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010110000000100101)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010110000000100110)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010110000000100111)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010110000000101000)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010110000000101001) && ({row_reg, col_reg}<18'b010110000000101100)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010110000000101100) && ({row_reg, col_reg}<18'b010110000000110001)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010110000000110001) && ({row_reg, col_reg}<18'b010110000000110011)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010110000000110011)) color_data = 12'b011111001110;
		if(({row_reg, col_reg}==18'b010110000000110100)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}==18'b010110000000110101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010110000000110110)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}==18'b010110000000110111)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==18'b010110000000111000)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010110000000111001)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010110000000111010)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010110000000111011)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010110000000111100)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}==18'b010110000000111101)) color_data = 12'b010110111101;
		if(({row_reg, col_reg}>=18'b010110000000111110) && ({row_reg, col_reg}<18'b010110000001000000)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}==18'b010110000001000000)) color_data = 12'b010010111011;
		if(({row_reg, col_reg}==18'b010110000001000001)) color_data = 12'b011011011101;
		if(({row_reg, col_reg}>=18'b010110000001000010) && ({row_reg, col_reg}<18'b010110000001000100)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010110000001000100) && ({row_reg, col_reg}<18'b010110000001000110)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010110000001000110) && ({row_reg, col_reg}<18'b010110000001001000)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010110000001001000)) color_data = 12'b100011111110;
		if(({row_reg, col_reg}==18'b010110000001001001)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010110000001001010)) color_data = 12'b011111111110;
		if(({row_reg, col_reg}>=18'b010110000001001011) && ({row_reg, col_reg}<18'b010110000001010001)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010110000001010001)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010110000001010010)) color_data = 12'b100011111110;
		if(({row_reg, col_reg}==18'b010110000001010011)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010110000001010100)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}==18'b010110000001010101)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}>=18'b010110000001010110) && ({row_reg, col_reg}<18'b010110000001011000)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010110000001011000)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b010110000001011001)) color_data = 12'b011011001110;
		if(({row_reg, col_reg}>=18'b010110000001011010) && ({row_reg, col_reg}<18'b010110000001011100)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010110000001011100)) color_data = 12'b100111111110;
		if(({row_reg, col_reg}==18'b010110000001011101)) color_data = 12'b101011101101;
		if(({row_reg, col_reg}>=18'b010110000001011110) && ({row_reg, col_reg}<18'b010110000001100000)) color_data = 12'b100110111011;
		if(({row_reg, col_reg}==18'b010110000001100000)) color_data = 12'b101010101000;
		if(({row_reg, col_reg}==18'b010110000001100001)) color_data = 12'b101010111001;
		if(({row_reg, col_reg}==18'b010110000001100010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010110000001100011) && ({row_reg, col_reg}<18'b010110000001100110)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==18'b010110000001100110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010110000001100111)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010110000001101000)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==18'b010110000001101001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010110000001101010)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==18'b010110000001101011)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010110000001101100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010110000001101101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010110000001101110) && ({row_reg, col_reg}<18'b010110000001110000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010110000001110000)) color_data = 12'b011001110101;
		if(({row_reg, col_reg}==18'b010110000001110001)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010110000001110010) && ({row_reg, col_reg}<18'b010110000001110101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010110000001110101)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b010110000001110110) && ({row_reg, col_reg}<18'b010110000001111000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010110000001111000)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}==18'b010110000001111001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010110000001111010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}>=18'b010110000001111011) && ({row_reg, col_reg}<18'b010110000001111101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010110000001111101)) color_data = 12'b101010111011;
		if(({row_reg, col_reg}==18'b010110000001111110)) color_data = 12'b100110101100;
		if(({row_reg, col_reg}==18'b010110000001111111)) color_data = 12'b011110001011;
		if(({row_reg, col_reg}>=18'b010110000010000000) && ({row_reg, col_reg}<18'b010110000010000010)) color_data = 12'b001101111010;
		if(({row_reg, col_reg}==18'b010110000010000010)) color_data = 12'b001110001011;
		if(({row_reg, col_reg}==18'b010110000010000011)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b010110000010000100)) color_data = 12'b011011011110;
		if(({row_reg, col_reg}>=18'b010110000010000101) && ({row_reg, col_reg}<18'b010110000010001000)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010110000010001000)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}==18'b010110000010001001)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b010110000010001010)) color_data = 12'b000101111011;
		if(({row_reg, col_reg}==18'b010110000010001011)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b010110000010001100)) color_data = 12'b000101111011;
		if(({row_reg, col_reg}==18'b010110000010001101)) color_data = 12'b010010101100;
		if(({row_reg, col_reg}==18'b010110000010001110)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010110000010001111)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}>=18'b010110000010010000) && ({row_reg, col_reg}<18'b010110000010010010)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010110000010010010)) color_data = 12'b010110111110;
		if(({row_reg, col_reg}==18'b010110000010010011)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}>=18'b010110000010010100) && ({row_reg, col_reg}<18'b010110000010010111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010110000010010111)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b010110000010011000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010110000010011001)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010110000010011010)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b010110000010011011)) color_data = 12'b001110011011;
		if(({row_reg, col_reg}==18'b010110000010011100)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010110000010011101)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010110000010011110) && ({row_reg, col_reg}<18'b010110000010100000)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010110000010100000) && ({row_reg, col_reg}<18'b010110000010100100)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010110000010100100) && ({row_reg, col_reg}<18'b010110000010100110)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010110000010100110)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010110000010100111) && ({row_reg, col_reg}<18'b010110000010101010)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010110000010101010)) color_data = 12'b010010101101;
		if(({row_reg, col_reg}==18'b010110000010101011)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b010110000010101100) && ({row_reg, col_reg}<18'b010110000010101110)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}>=18'b010110000010101110) && ({row_reg, col_reg}<18'b010110000010110000)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b010110000010110000)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b010110000010110001)) color_data = 12'b000101111100;
		if(({row_reg, col_reg}>=18'b010110000010110010) && ({row_reg, col_reg}<18'b010110000010110100)) color_data = 12'b001010001101;
		if(({row_reg, col_reg}==18'b010110000010110100)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b010110000010110101)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010110000010110110)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010110000010110111)) color_data = 12'b010001111011;
		if(({row_reg, col_reg}==18'b010110000010111000)) color_data = 12'b010001111010;
		if(({row_reg, col_reg}==18'b010110000010111001)) color_data = 12'b010101111000;
		if(({row_reg, col_reg}==18'b010110000010111010)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}>=18'b010110000010111011) && ({row_reg, col_reg}<18'b010110000010111110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010110000010111110)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}==18'b010110000010111111)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}>=18'b010110000011000000) && ({row_reg, col_reg}<18'b010110000011000010)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010110000011000010) && ({row_reg, col_reg}<18'b010110000011001011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010110000011001011)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010110000011001100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010110000011001101)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}>=18'b010110000011001110) && ({row_reg, col_reg}<18'b010110000011010000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010110000011010000)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==18'b010110000011010001)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}==18'b010110000011010010)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010110000011010011) && ({row_reg, col_reg}<18'b010110000011010101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010110000011010101) && ({row_reg, col_reg}<18'b010110000011100000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010110000011100000) && ({row_reg, col_reg}<18'b010110000011100010)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010110000011100010) && ({row_reg, col_reg}<18'b010110000011101001)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010110000011101001)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010110000011101010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010110000011101011) && ({row_reg, col_reg}<18'b010110000011101110)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}==18'b010110000011101110)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==18'b010110000011101111)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}>=18'b010110000011110000) && ({row_reg, col_reg}<18'b010110000011110010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010110000011110010)) color_data = 12'b010101100111;
		if(({row_reg, col_reg}==18'b010110000011110011)) color_data = 12'b011001111000;
		if(({row_reg, col_reg}==18'b010110000011110100)) color_data = 12'b010110001000;
		if(({row_reg, col_reg}==18'b010110000011110101)) color_data = 12'b001101110111;
		if(({row_reg, col_reg}==18'b010110000011110110)) color_data = 12'b011010111011;
		if(({row_reg, col_reg}==18'b010110000011110111)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010110000011111000)) color_data = 12'b100111111110;
		if(({row_reg, col_reg}==18'b010110000011111001)) color_data = 12'b100011111110;
		if(({row_reg, col_reg}==18'b010110000011111010)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010110000011111011)) color_data = 12'b010110111101;
		if(({row_reg, col_reg}==18'b010110000011111100)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b010110000011111101) && ({row_reg, col_reg}<18'b010110000011111111)) color_data = 12'b001010001101;
		if(({row_reg, col_reg}==18'b010110000011111111)) color_data = 12'b001010011101;
		if(({row_reg, col_reg}==18'b010110000100000000)) color_data = 12'b100011101110;
		if(({row_reg, col_reg}>=18'b010110000100000001) && ({row_reg, col_reg}<18'b010110000100000011)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010110000100000011) && ({row_reg, col_reg}<18'b010110000100000110)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010110000100000110)) color_data = 12'b011111111111;
		if(({row_reg, col_reg}==18'b010110000100000111)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010110000100001000)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010110000100001001)) color_data = 12'b100011011110;
		if(({row_reg, col_reg}==18'b010110000100001010)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}==18'b010110000100001011)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==18'b010110000100001100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010110000100001101) && ({row_reg, col_reg}<18'b010110000100001111)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b010110000100001111)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}==18'b010110000100010000)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b010110000100010001) && ({row_reg, col_reg}<18'b010110001000000010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010110001000000010)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b010110001000000011)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}==18'b010110001000000100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010110001000000101) && ({row_reg, col_reg}<18'b010110001000001000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010110001000001000) && ({row_reg, col_reg}<18'b010110001000001111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010110001000001111)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010110001000010000) && ({row_reg, col_reg}<18'b010110001000010010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010110001000010010)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}>=18'b010110001000010011) && ({row_reg, col_reg}<18'b010110001000010101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010110001000010101) && ({row_reg, col_reg}<18'b010110001000100000)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b010110001000100000)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010110001000100001)) color_data = 12'b011111101111;
		if(({row_reg, col_reg}>=18'b010110001000100010) && ({row_reg, col_reg}<18'b010110001000100100)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010110001000100100)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010110001000100101)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010110001000100110)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010110001000100111)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010110001000101000) && ({row_reg, col_reg}<18'b010110001000101101)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}>=18'b010110001000101101) && ({row_reg, col_reg}<18'b010110001000110001)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010110001000110001)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010110001000110010)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b010110001000110011)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==18'b010110001000110100)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}==18'b010110001000110101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010110001000110110)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==18'b010110001000110111)) color_data = 12'b011111001111;
		if(({row_reg, col_reg}>=18'b010110001000111000) && ({row_reg, col_reg}<18'b010110001000111010)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}>=18'b010110001000111010) && ({row_reg, col_reg}<18'b010110001000111100)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010110001000111100)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}==18'b010110001000111101)) color_data = 12'b011011001110;
		if(({row_reg, col_reg}==18'b010110001000111110)) color_data = 12'b010110111101;
		if(({row_reg, col_reg}==18'b010110001000111111)) color_data = 12'b010110101100;
		if(({row_reg, col_reg}==18'b010110001001000000)) color_data = 12'b010111001100;
		if(({row_reg, col_reg}==18'b010110001001000001)) color_data = 12'b011111011110;
		if(({row_reg, col_reg}==18'b010110001001000010)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010110001001000011)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010110001001000100)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010110001001000101) && ({row_reg, col_reg}<18'b010110001001001100)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010110001001001100)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}>=18'b010110001001001101) && ({row_reg, col_reg}<18'b010110001001010001)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010110001001010001) && ({row_reg, col_reg}<18'b010110001001010011)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010110001001010011)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010110001001010100)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}>=18'b010110001001010101) && ({row_reg, col_reg}<18'b010110001001011000)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b010110001001011000)) color_data = 12'b001110011100;
		if(({row_reg, col_reg}==18'b010110001001011001)) color_data = 12'b010111001110;
		if(({row_reg, col_reg}>=18'b010110001001011010) && ({row_reg, col_reg}<18'b010110001001011100)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010110001001011100)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b010110001001011101)) color_data = 12'b100111011101;
		if(({row_reg, col_reg}==18'b010110001001011110)) color_data = 12'b100111001100;
		if(({row_reg, col_reg}==18'b010110001001011111)) color_data = 12'b100110111011;
		if(({row_reg, col_reg}==18'b010110001001100000)) color_data = 12'b101010111001;
		if(({row_reg, col_reg}==18'b010110001001100001)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==18'b010110001001100010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010110001001100011)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==18'b010110001001100100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010110001001100101)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==18'b010110001001100110)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}>=18'b010110001001100111) && ({row_reg, col_reg}<18'b010110001001101001)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}>=18'b010110001001101001) && ({row_reg, col_reg}<18'b010110001001101100)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010110001001101100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010110001001101101) && ({row_reg, col_reg}<18'b010110001001110000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010110001001110000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010110001001110001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010110001001110010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010110001001110011)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}==18'b010110001001110100)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010110001001110101)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010110001001110110)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010110001001110111)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010110001001111000)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010110001001111001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010110001001111010)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010110001001111011)) color_data = 12'b101110111010;
		if(({row_reg, col_reg}==18'b010110001001111100)) color_data = 12'b101010111010;
		if(({row_reg, col_reg}==18'b010110001001111101)) color_data = 12'b101010111011;
		if(({row_reg, col_reg}==18'b010110001001111110)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b010110001001111111)) color_data = 12'b011110001010;
		if(({row_reg, col_reg}==18'b010110001010000000)) color_data = 12'b010010001011;
		if(({row_reg, col_reg}==18'b010110001010000001)) color_data = 12'b001110001011;
		if(({row_reg, col_reg}==18'b010110001010000010)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b010110001010000011)) color_data = 12'b001010011011;
		if(({row_reg, col_reg}==18'b010110001010000100)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}>=18'b010110001010000101) && ({row_reg, col_reg}<18'b010110001010001000)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010110001010001000)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}==18'b010110001010001001)) color_data = 12'b001110011100;
		if(({row_reg, col_reg}==18'b010110001010001010)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b010110001010001011)) color_data = 12'b000110001011;
		if(({row_reg, col_reg}==18'b010110001010001100)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b010110001010001101)) color_data = 12'b010110111101;
		if(({row_reg, col_reg}==18'b010110001010001110)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010110001010001111)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b010110001010010000)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010110001010010001)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010110001010010010)) color_data = 12'b010110101101;
		if(({row_reg, col_reg}==18'b010110001010010011)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b010110001010010100) && ({row_reg, col_reg}<18'b010110001010011000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010110001010011000)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010110001010011001)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010110001010011010)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010110001010011011)) color_data = 12'b001110011011;
		if(({row_reg, col_reg}==18'b010110001010011100)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}>=18'b010110001010011101) && ({row_reg, col_reg}<18'b010110001010011111)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010110001010011111) && ({row_reg, col_reg}<18'b010110001010100001)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010110001010100001)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010110001010100010) && ({row_reg, col_reg}<18'b010110001010101001)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010110001010101001)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010110001010101010)) color_data = 12'b010111001110;
		if(({row_reg, col_reg}==18'b010110001010101011)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b010110001010101100)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b010110001010101101)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b010110001010101110)) color_data = 12'b001010001010;
		if(({row_reg, col_reg}==18'b010110001010101111)) color_data = 12'b001010011011;
		if(({row_reg, col_reg}==18'b010110001010110000)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b010110001010110001)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}>=18'b010110001010110010) && ({row_reg, col_reg}<18'b010110001010110110)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b010110001010110110)) color_data = 12'b001110001011;
		if(({row_reg, col_reg}==18'b010110001010110111)) color_data = 12'b001101111010;
		if(({row_reg, col_reg}==18'b010110001010111000)) color_data = 12'b010001111001;
		if(({row_reg, col_reg}==18'b010110001010111001)) color_data = 12'b010101111000;
		if(({row_reg, col_reg}==18'b010110001010111010)) color_data = 12'b010101110111;
		if(({row_reg, col_reg}==18'b010110001010111011)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==18'b010110001010111100)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}>=18'b010110001010111101) && ({row_reg, col_reg}<18'b010110001011000000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010110001011000000)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010110001011000001) && ({row_reg, col_reg}<18'b010110001011000011)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010110001011000011) && ({row_reg, col_reg}<18'b010110001011100000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010110001011100000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010110001011100001)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010110001011100010) && ({row_reg, col_reg}<18'b010110001011101010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010110001011101010)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}==18'b010110001011101011)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==18'b010110001011101100)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}==18'b010110001011101101)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==18'b010110001011101110)) color_data = 12'b011001111000;
		if(({row_reg, col_reg}==18'b010110001011101111)) color_data = 12'b011001101000;
		if(({row_reg, col_reg}==18'b010110001011110000)) color_data = 12'b010101100111;
		if(({row_reg, col_reg}==18'b010110001011110001)) color_data = 12'b010101111000;
		if(({row_reg, col_reg}==18'b010110001011110010)) color_data = 12'b011010001001;
		if(({row_reg, col_reg}==18'b010110001011110011)) color_data = 12'b010110001000;
		if(({row_reg, col_reg}==18'b010110001011110100)) color_data = 12'b010001111000;
		if(({row_reg, col_reg}==18'b010110001011110101)) color_data = 12'b001101111000;
		if(({row_reg, col_reg}==18'b010110001011110110)) color_data = 12'b010110101010;
		if(({row_reg, col_reg}==18'b010110001011110111)) color_data = 12'b100111101110;
		if(({row_reg, col_reg}==18'b010110001011111000)) color_data = 12'b100111111110;
		if(({row_reg, col_reg}>=18'b010110001011111001) && ({row_reg, col_reg}<18'b010110001011111011)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010110001011111011)) color_data = 12'b010010101101;
		if(({row_reg, col_reg}==18'b010110001011111100)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010110001011111101)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010110001011111110)) color_data = 12'b000101111100;
		if(({row_reg, col_reg}==18'b010110001011111111)) color_data = 12'b001010001101;
		if(({row_reg, col_reg}==18'b010110001100000000)) color_data = 12'b011111101110;
		if(({row_reg, col_reg}>=18'b010110001100000001) && ({row_reg, col_reg}<18'b010110001100000100)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010110001100000100) && ({row_reg, col_reg}<18'b010110001100001000)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010110001100001000)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010110001100001001)) color_data = 12'b011111011110;
		if(({row_reg, col_reg}==18'b010110001100001010)) color_data = 12'b010110101101;
		if(({row_reg, col_reg}>=18'b010110001100001011) && ({row_reg, col_reg}<18'b010110001100001110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010110001100001110)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b010110001100001111)) color_data = 12'b011110101111;

		if(({row_reg, col_reg}>=18'b010110001100010000) && ({row_reg, col_reg}<18'b010110010000001010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010110010000001010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010110010000001011) && ({row_reg, col_reg}<18'b010110010000001111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010110010000001111)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b010110010000010000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010110010000010001)) color_data = 12'b010110011101;
		if(({row_reg, col_reg}>=18'b010110010000010010) && ({row_reg, col_reg}<18'b010110010000010100)) color_data = 12'b010010001100;
		if(({row_reg, col_reg}>=18'b010110010000010100) && ({row_reg, col_reg}<18'b010110010000010110)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}>=18'b010110010000010110) && ({row_reg, col_reg}<18'b010110010000011000)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}>=18'b010110010000011000) && ({row_reg, col_reg}<18'b010110010000011010)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010110010000011010)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}>=18'b010110010000011011) && ({row_reg, col_reg}<18'b010110010000011101)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}==18'b010110010000011101)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b010110010000011110)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010110010000011111)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010110010000100000)) color_data = 12'b001110011101;
		if(({row_reg, col_reg}==18'b010110010000100001)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}>=18'b010110010000100010) && ({row_reg, col_reg}<18'b010110010000100100)) color_data = 12'b001110011101;
		if(({row_reg, col_reg}>=18'b010110010000100100) && ({row_reg, col_reg}<18'b010110010000110001)) color_data = 12'b001110011100;
		if(({row_reg, col_reg}>=18'b010110010000110001) && ({row_reg, col_reg}<18'b010110010000110011)) color_data = 12'b010010011100;
		if(({row_reg, col_reg}==18'b010110010000110011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010110010000110100)) color_data = 12'b010110101101;
		if(({row_reg, col_reg}==18'b010110010000110101)) color_data = 12'b011110111111;
		if(({row_reg, col_reg}==18'b010110010000110110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010110010000110111)) color_data = 12'b010110101101;
		if(({row_reg, col_reg}==18'b010110010000111000)) color_data = 12'b010010011101;
		if(({row_reg, col_reg}>=18'b010110010000111001) && ({row_reg, col_reg}<18'b010110010000111011)) color_data = 12'b001110011100;
		if(({row_reg, col_reg}==18'b010110010000111011)) color_data = 12'b001110011011;
		if(({row_reg, col_reg}==18'b010110010000111100)) color_data = 12'b010110111101;
		if(({row_reg, col_reg}>=18'b010110010000111101) && ({row_reg, col_reg}<18'b010110010001000000)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010110010001000000)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010110010001000001)) color_data = 12'b011111101110;
		if(({row_reg, col_reg}>=18'b010110010001000010) && ({row_reg, col_reg}<18'b010110010001000100)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010110010001000100)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010110010001000101)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010110010001000110)) color_data = 12'b010110111101;
		if(({row_reg, col_reg}==18'b010110010001000111)) color_data = 12'b001110011100;
		if(({row_reg, col_reg}==18'b010110010001001000)) color_data = 12'b001010011011;
		if(({row_reg, col_reg}==18'b010110010001001001)) color_data = 12'b001010011100;
		if(({row_reg, col_reg}>=18'b010110010001001010) && ({row_reg, col_reg}<18'b010110010001010000)) color_data = 12'b001110011100;
		if(({row_reg, col_reg}==18'b010110010001010000)) color_data = 12'b001110011101;
		if(({row_reg, col_reg}==18'b010110010001010001)) color_data = 12'b001110011100;
		if(({row_reg, col_reg}==18'b010110010001010010)) color_data = 12'b010010011100;
		if(({row_reg, col_reg}==18'b010110010001010011)) color_data = 12'b010010011011;
		if(({row_reg, col_reg}==18'b010110010001010100)) color_data = 12'b010110111101;
		if(({row_reg, col_reg}==18'b010110010001010101)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}>=18'b010110010001010110) && ({row_reg, col_reg}<18'b010110010001011000)) color_data = 12'b100011011111;
		if(({row_reg, col_reg}==18'b010110010001011000)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}==18'b010110010001011001)) color_data = 12'b010010111101;
		if(({row_reg, col_reg}>=18'b010110010001011010) && ({row_reg, col_reg}<18'b010110010001011100)) color_data = 12'b001110011011;
		if(({row_reg, col_reg}==18'b010110010001011100)) color_data = 12'b010010011011;
		if(({row_reg, col_reg}==18'b010110010001011101)) color_data = 12'b011010011011;
		if(({row_reg, col_reg}>=18'b010110010001011110) && ({row_reg, col_reg}<18'b010110010001100000)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}>=18'b010110010001100000) && ({row_reg, col_reg}<18'b010110010001100010)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010110010001100010)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010110010001100011) && ({row_reg, col_reg}<18'b010110010001100110)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}>=18'b010110010001100110) && ({row_reg, col_reg}<18'b010110010001101000)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010110010001101000)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010110010001101001)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}==18'b010110010001101010)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==18'b010110010001101011)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010110010001101100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010110010001101101)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==18'b010110010001101110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010110010001101111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010110010001110000)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010110010001110001) && ({row_reg, col_reg}<18'b010110010001110100)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}==18'b010110010001110100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010110010001110101)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010110010001110110) && ({row_reg, col_reg}<18'b010110010001111010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010110010001111010)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}==18'b010110010001111011)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==18'b010110010001111100)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010110010001111101)) color_data = 12'b101010111010;
		if(({row_reg, col_reg}==18'b010110010001111110)) color_data = 12'b100110111011;
		if(({row_reg, col_reg}==18'b010110010001111111)) color_data = 12'b100110111100;
		if(({row_reg, col_reg}==18'b010110010010000000)) color_data = 12'b100011001111;
		if(({row_reg, col_reg}==18'b010110010010000001)) color_data = 12'b100011011111;
		if(({row_reg, col_reg}==18'b010110010010000010)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010110010010000011)) color_data = 12'b011111101111;
		if(({row_reg, col_reg}>=18'b010110010010000100) && ({row_reg, col_reg}<18'b010110010010001000)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010110010010001000)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010110010010001001)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}==18'b010110010010001010)) color_data = 12'b011111101111;
		if(({row_reg, col_reg}==18'b010110010010001011)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010110010010001100)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}==18'b010110010010001101)) color_data = 12'b010111001110;
		if(({row_reg, col_reg}==18'b010110010010001110)) color_data = 12'b010010101101;
		if(({row_reg, col_reg}==18'b010110010010001111)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b010110010010010000)) color_data = 12'b001110011100;
		if(({row_reg, col_reg}==18'b010110010010010001)) color_data = 12'b010010101101;
		if(({row_reg, col_reg}==18'b010110010010010010)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}>=18'b010110010010010011) && ({row_reg, col_reg}<18'b010110010010010101)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010110010010010101)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010110010010010110)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b010110010010010111) && ({row_reg, col_reg}<18'b010110010010011001)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010110010010011001)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010110010010011010)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010110010010011011)) color_data = 12'b001110011100;
		if(({row_reg, col_reg}==18'b010110010010011100)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010110010010011101)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010110010010011110) && ({row_reg, col_reg}<18'b010110010010100001)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010110010010100001)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010110010010100010) && ({row_reg, col_reg}<18'b010110010010101010)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010110010010101010)) color_data = 12'b011111101111;
		if(({row_reg, col_reg}==18'b010110010010101011)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}==18'b010110010010101100)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}>=18'b010110010010101101) && ({row_reg, col_reg}<18'b010110010010101111)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}==18'b010110010010101111)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010110010010110000)) color_data = 12'b011111101111;
		if(({row_reg, col_reg}==18'b010110010010110001)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}>=18'b010110010010110010) && ({row_reg, col_reg}<18'b010110010010110100)) color_data = 12'b011111101111;
		if(({row_reg, col_reg}>=18'b010110010010110100) && ({row_reg, col_reg}<18'b010110010010110110)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}>=18'b010110010010110110) && ({row_reg, col_reg}<18'b010110010010111000)) color_data = 12'b100011011111;
		if(({row_reg, col_reg}==18'b010110010010111000)) color_data = 12'b100011011110;
		if(({row_reg, col_reg}==18'b010110010010111001)) color_data = 12'b100111011110;
		if(({row_reg, col_reg}==18'b010110010010111010)) color_data = 12'b101011011110;
		if(({row_reg, col_reg}==18'b010110010010111011)) color_data = 12'b101111011101;
		if(({row_reg, col_reg}==18'b010110010010111100)) color_data = 12'b101011001100;
		if(({row_reg, col_reg}==18'b010110010010111101)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}==18'b010110010010111110)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}==18'b010110010010111111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010110010011000000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010110010011000001)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010110010011000010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010110010011000011)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==18'b010110010011000100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010110010011000101) && ({row_reg, col_reg}<18'b010110010011000111)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010110010011000111) && ({row_reg, col_reg}<18'b010110010011010000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010110010011010000) && ({row_reg, col_reg}<18'b010110010011010110)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010110010011010110) && ({row_reg, col_reg}<18'b010110010011100000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010110010011100000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010110010011100001)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010110010011100010) && ({row_reg, col_reg}<18'b010110010011101001)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010110010011101001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010110010011101010)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}==18'b010110010011101011)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==18'b010110010011101100)) color_data = 12'b010101110111;
		if(({row_reg, col_reg}==18'b010110010011101101)) color_data = 12'b010101111000;
		if(({row_reg, col_reg}>=18'b010110010011101110) && ({row_reg, col_reg}<18'b010110010011110001)) color_data = 12'b010101111001;
		if(({row_reg, col_reg}==18'b010110010011110001)) color_data = 12'b011110011011;
		if(({row_reg, col_reg}==18'b010110010011110010)) color_data = 12'b100111001101;
		if(({row_reg, col_reg}>=18'b010110010011110011) && ({row_reg, col_reg}<18'b010110010011110101)) color_data = 12'b100111011101;
		if(({row_reg, col_reg}==18'b010110010011110101)) color_data = 12'b100011011101;
		if(({row_reg, col_reg}==18'b010110010011110110)) color_data = 12'b100111101110;
		if(({row_reg, col_reg}==18'b010110010011110111)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010110010011111000)) color_data = 12'b100011111110;
		if(({row_reg, col_reg}==18'b010110010011111001)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010110010011111010)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010110010011111011)) color_data = 12'b010010101101;
		if(({row_reg, col_reg}>=18'b010110010011111100) && ({row_reg, col_reg}<18'b010110010011111110)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010110010011111110)) color_data = 12'b001010001101;
		if(({row_reg, col_reg}==18'b010110010011111111)) color_data = 12'b001110011101;
		if(({row_reg, col_reg}==18'b010110010100000000)) color_data = 12'b011111101110;
		if(({row_reg, col_reg}>=18'b010110010100000001) && ({row_reg, col_reg}<18'b010110010100000110)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010110010100000110)) color_data = 12'b100011111110;
		if(({row_reg, col_reg}>=18'b010110010100000111) && ({row_reg, col_reg}<18'b010110010100001001)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010110010100001001)) color_data = 12'b011011001110;
		if(({row_reg, col_reg}==18'b010110010100001010)) color_data = 12'b001110001011;
		if(({row_reg, col_reg}>=18'b010110010100001011) && ({row_reg, col_reg}<18'b010110010100001101)) color_data = 12'b010010001100;
		if(({row_reg, col_reg}==18'b010110010100001101)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}==18'b010110010100001110)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==18'b010110010100001111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010110010100010000)) color_data = 12'b011110111111;
		if(({row_reg, col_reg}==18'b010110010100010001)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b010110010100010010) && ({row_reg, col_reg}<18'b010110011000001010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010110011000001010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010110011000001011) && ({row_reg, col_reg}<18'b010110011000010000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010110011000010000)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b010110011000010001)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==18'b010110011000010010)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}>=18'b010110011000010011) && ({row_reg, col_reg}<18'b010110011000010101)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}>=18'b010110011000010101) && ({row_reg, col_reg}<18'b010110011000100000)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010110011000100000)) color_data = 12'b001010001101;
		if(({row_reg, col_reg}>=18'b010110011000100001) && ({row_reg, col_reg}<18'b010110011000100110)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010110011000100110) && ({row_reg, col_reg}<18'b010110011000101100)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b010110011000101100) && ({row_reg, col_reg}<18'b010110011000101110)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010110011000101110) && ({row_reg, col_reg}<18'b010110011000110010)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010110011000110010)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010110011000110011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010110011000110100)) color_data = 12'b011110111111;
		if(({row_reg, col_reg}==18'b010110011000110101)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b010110011000110110)) color_data = 12'b011010011110;
		if(({row_reg, col_reg}==18'b010110011000110111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010110011000111000)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}>=18'b010110011000111001) && ({row_reg, col_reg}<18'b010110011000111011)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b010110011000111011)) color_data = 12'b000101111010;
		if(({row_reg, col_reg}==18'b010110011000111100)) color_data = 12'b010010101100;
		if(({row_reg, col_reg}>=18'b010110011000111101) && ({row_reg, col_reg}<18'b010110011000111111)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010110011000111111) && ({row_reg, col_reg}<18'b010110011001000011)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010110011001000011) && ({row_reg, col_reg}<18'b010110011001000101)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010110011001000101)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010110011001000110)) color_data = 12'b010010101100;
		if(({row_reg, col_reg}==18'b010110011001000111)) color_data = 12'b000101111010;
		if(({row_reg, col_reg}==18'b010110011001001000)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b010110011001001001)) color_data = 12'b000101111100;
		if(({row_reg, col_reg}>=18'b010110011001001010) && ({row_reg, col_reg}<18'b010110011001001100)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010110011001001100)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}>=18'b010110011001001101) && ({row_reg, col_reg}<18'b010110011001010000)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010110011001010000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010110011001010001) && ({row_reg, col_reg}<18'b010110011001010011)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010110011001010011)) color_data = 12'b001001111010;
		if(({row_reg, col_reg}==18'b010110011001010100)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}>=18'b010110011001010101) && ({row_reg, col_reg}<18'b010110011001011001)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010110011001011001)) color_data = 12'b010010101100;
		if(({row_reg, col_reg}==18'b010110011001011010)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b010110011001011011)) color_data = 12'b000101111010;
		if(({row_reg, col_reg}==18'b010110011001011100)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b010110011001011101)) color_data = 12'b010001111010;
		if(({row_reg, col_reg}==18'b010110011001011110)) color_data = 12'b100010011100;
		if(({row_reg, col_reg}==18'b010110011001011111)) color_data = 12'b100010011011;
		if(({row_reg, col_reg}==18'b010110011001100000)) color_data = 12'b101010011010;
		if(({row_reg, col_reg}==18'b010110011001100001)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010110011001100010) && ({row_reg, col_reg}<18'b010110011001100101)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010110011001100101)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010110011001100110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010110011001100111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010110011001101000)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}>=18'b010110011001101001) && ({row_reg, col_reg}<18'b010110011001101011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010110011001101011)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==18'b010110011001101100)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}==18'b010110011001101101)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}>=18'b010110011001101110) && ({row_reg, col_reg}<18'b010110011001110000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010110011001110000)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010110011001110001) && ({row_reg, col_reg}<18'b010110011001110100)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}==18'b010110011001110100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010110011001110101)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==18'b010110011001110110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010110011001110111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010110011001111000)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==18'b010110011001111001)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010110011001111010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010110011001111011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010110011001111100)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010110011001111101)) color_data = 12'b101010111010;
		if(({row_reg, col_reg}==18'b010110011001111110)) color_data = 12'b100110111011;
		if(({row_reg, col_reg}==18'b010110011001111111)) color_data = 12'b101011001101;
		if(({row_reg, col_reg}>=18'b010110011010000000) && ({row_reg, col_reg}<18'b010110011010000010)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}==18'b010110011010000010)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010110011010000011) && ({row_reg, col_reg}<18'b010110011010001000)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010110011010001000)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010110011010001001)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010110011010001010) && ({row_reg, col_reg}<18'b010110011010001100)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010110011010001100)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010110011010001101)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}==18'b010110011010001110)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b010110011010001111)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}>=18'b010110011010010000) && ({row_reg, col_reg}<18'b010110011010010011)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010110011010010011)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010110011010010100) && ({row_reg, col_reg}<18'b010110011010010110)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b010110011010010110)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010110011010010111) && ({row_reg, col_reg}<18'b010110011010011010)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010110011010011010)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010110011010011011)) color_data = 12'b001110011100;
		if(({row_reg, col_reg}==18'b010110011010011100)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010110011010011101)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010110011010011110) && ({row_reg, col_reg}<18'b010110011010100000)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010110011010100000)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010110011010100001) && ({row_reg, col_reg}<18'b010110011010101011)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010110011010101011) && ({row_reg, col_reg}<18'b010110011010111001)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010110011010111001)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b010110011010111010)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}==18'b010110011010111011)) color_data = 12'b101111101111;
		if(({row_reg, col_reg}==18'b010110011010111100)) color_data = 12'b110011101111;
		if(({row_reg, col_reg}==18'b010110011010111101)) color_data = 12'b011110011001;
		if(({row_reg, col_reg}>=18'b010110011010111110) && ({row_reg, col_reg}<18'b010110011011000000)) color_data = 12'b010101110110;
		if(({row_reg, col_reg}==18'b010110011011000000)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}>=18'b010110011011000001) && ({row_reg, col_reg}<18'b010110011011000011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010110011011000011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010110011011000100) && ({row_reg, col_reg}<18'b010110011011000111)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==18'b010110011011000111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010110011011001000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010110011011001001) && ({row_reg, col_reg}<18'b010110011011001101)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010110011011001101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010110011011001110) && ({row_reg, col_reg}<18'b010110011011010111)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010110011011010111) && ({row_reg, col_reg}<18'b010110011011011110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010110011011011110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010110011011011111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010110011011100000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010110011011100001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010110011011100010) && ({row_reg, col_reg}<18'b010110011011100101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010110011011100101) && ({row_reg, col_reg}<18'b010110011011100111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010110011011100111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010110011011101000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010110011011101001) && ({row_reg, col_reg}<18'b010110011011101011)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}==18'b010110011011101011)) color_data = 12'b010101110111;
		if(({row_reg, col_reg}==18'b010110011011101100)) color_data = 12'b010101111000;
		if(({row_reg, col_reg}==18'b010110011011101101)) color_data = 12'b010001111001;
		if(({row_reg, col_reg}>=18'b010110011011101110) && ({row_reg, col_reg}<18'b010110011011110000)) color_data = 12'b010001111010;
		if(({row_reg, col_reg}==18'b010110011011110000)) color_data = 12'b001101101010;
		if(({row_reg, col_reg}==18'b010110011011110001)) color_data = 12'b010110011100;
		if(({row_reg, col_reg}==18'b010110011011110010)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}==18'b010110011011110011)) color_data = 12'b101011111110;
		if(({row_reg, col_reg}==18'b010110011011110100)) color_data = 12'b100111111110;
		if(({row_reg, col_reg}==18'b010110011011110101)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010110011011110110)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010110011011110111)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010110011011111000)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010110011011111001) && ({row_reg, col_reg}<18'b010110011011111011)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010110011011111011)) color_data = 12'b010010101110;
		if(({row_reg, col_reg}>=18'b010110011011111100) && ({row_reg, col_reg}<18'b010110011011111110)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010110011011111110)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010110011011111111)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b010110011100000000)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}>=18'b010110011100000001) && ({row_reg, col_reg}<18'b010110011100000101)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010110011100000101)) color_data = 12'b100011111110;
		if(({row_reg, col_reg}==18'b010110011100000110)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010110011100000111)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010110011100001000)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010110011100001001)) color_data = 12'b011011001110;
		if(({row_reg, col_reg}==18'b010110011100001010)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}>=18'b010110011100001011) && ({row_reg, col_reg}<18'b010110011100001110)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010110011100001110)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==18'b010110011100001111)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b010110011100010000)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b010110011100010001) && ({row_reg, col_reg}<18'b010110100000010000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010110100000010000)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b010110100000010001)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==18'b010110100000010010)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010110100000010011)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}>=18'b010110100000010100) && ({row_reg, col_reg}<18'b010110100000010111)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010110100000010111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010110100000011000) && ({row_reg, col_reg}<18'b010110100000011011)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b010110100000011011) && ({row_reg, col_reg}<18'b010110100000011110)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b010110100000011110) && ({row_reg, col_reg}<18'b010110100000100000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010110100000100000)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b010110100000100001)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}>=18'b010110100000100010) && ({row_reg, col_reg}<18'b010110100000100111)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}>=18'b010110100000100111) && ({row_reg, col_reg}<18'b010110100000101001)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010110100000101001) && ({row_reg, col_reg}<18'b010110100000101111)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010110100000101111)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}>=18'b010110100000110000) && ({row_reg, col_reg}<18'b010110100000110010)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010110100000110010)) color_data = 12'b010001111101;
		if(({row_reg, col_reg}==18'b010110100000110011)) color_data = 12'b010110001101;
		if(({row_reg, col_reg}>=18'b010110100000110100) && ({row_reg, col_reg}<18'b010110100000110110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010110100000110110)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b010110100000110111)) color_data = 12'b011010111111;
		if(({row_reg, col_reg}==18'b010110100000111000)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010110100000111001)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010110100000111010)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b010110100000111011)) color_data = 12'b001010001010;
		if(({row_reg, col_reg}==18'b010110100000111100)) color_data = 12'b010110111101;
		if(({row_reg, col_reg}>=18'b010110100000111101) && ({row_reg, col_reg}<18'b010110100001000000)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010110100001000000) && ({row_reg, col_reg}<18'b010110100001000010)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010110100001000010)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010110100001000011) && ({row_reg, col_reg}<18'b010110100001000110)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010110100001000110)) color_data = 12'b010010101101;
		if(({row_reg, col_reg}==18'b010110100001000111)) color_data = 12'b000101111011;
		if(({row_reg, col_reg}==18'b010110100001001000)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b010110100001001001)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010110100001001010)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}>=18'b010110100001001011) && ({row_reg, col_reg}<18'b010110100001010000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010110100001010000)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b010110100001010001)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010110100001010010)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010110100001010011)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b010110100001010100)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==18'b010110100001010101)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}>=18'b010110100001010110) && ({row_reg, col_reg}<18'b010110100001011000)) color_data = 12'b100011101110;
		if(({row_reg, col_reg}==18'b010110100001011000)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010110100001011001)) color_data = 12'b010010101100;
		if(({row_reg, col_reg}==18'b010110100001011010)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b010110100001011011)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b010110100001011100)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}==18'b010110100001011101)) color_data = 12'b010001111011;
		if(({row_reg, col_reg}==18'b010110100001011110)) color_data = 12'b100010101100;
		if(({row_reg, col_reg}==18'b010110100001011111)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}>=18'b010110100001100000) && ({row_reg, col_reg}<18'b010110100001100010)) color_data = 12'b101010011001;
		if(({row_reg, col_reg}==18'b010110100001100010)) color_data = 12'b101010011000;
		if(({row_reg, col_reg}>=18'b010110100001100011) && ({row_reg, col_reg}<18'b010110100001100110)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010110100001100110)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010110100001100111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010110100001101000)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}==18'b010110100001101001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010110100001101010) && ({row_reg, col_reg}<18'b010110100001101100)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}==18'b010110100001101100)) color_data = 12'b011101110101;
		if(({row_reg, col_reg}==18'b010110100001101101)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}>=18'b010110100001101110) && ({row_reg, col_reg}<18'b010110100001110000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010110100001110000)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010110100001110001) && ({row_reg, col_reg}<18'b010110100001110011)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}>=18'b010110100001110011) && ({row_reg, col_reg}<18'b010110100001110101)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010110100001110101)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}>=18'b010110100001110110) && ({row_reg, col_reg}<18'b010110100001111000)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}>=18'b010110100001111000) && ({row_reg, col_reg}<18'b010110100001111010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010110100001111010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010110100001111011)) color_data = 12'b101110101010;
		if(({row_reg, col_reg}==18'b010110100001111100)) color_data = 12'b101010111011;
		if(({row_reg, col_reg}>=18'b010110100001111101) && ({row_reg, col_reg}<18'b010110100001111111)) color_data = 12'b100110111011;
		if(({row_reg, col_reg}==18'b010110100001111111)) color_data = 12'b101011001101;
		if(({row_reg, col_reg}==18'b010110100010000000)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b010110100010000001)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010110100010000010) && ({row_reg, col_reg}<18'b010110100010001000)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010110100010001000) && ({row_reg, col_reg}<18'b010110100010001011)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010110100010001011)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010110100010001100)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010110100010001101)) color_data = 12'b011011011111;
		if(({row_reg, col_reg}>=18'b010110100010001110) && ({row_reg, col_reg}<18'b010110100010010000)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b010110100010010000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010110100010010001) && ({row_reg, col_reg}<18'b010110100010010011)) color_data = 12'b001010001101;
		if(({row_reg, col_reg}>=18'b010110100010010011) && ({row_reg, col_reg}<18'b010110100010010101)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010110100010010101)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010110100010010110)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010110100010010111) && ({row_reg, col_reg}<18'b010110100010011010)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010110100010011010)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010110100010011011)) color_data = 12'b001110011100;
		if(({row_reg, col_reg}==18'b010110100010011100)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010110100010011101)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010110100010011110) && ({row_reg, col_reg}<18'b010110100010100000)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010110100010100000)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010110100010100001) && ({row_reg, col_reg}<18'b010110100010100100)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010110100010100100)) color_data = 12'b100011111110;
		if(({row_reg, col_reg}>=18'b010110100010100101) && ({row_reg, col_reg}<18'b010110100010101011)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010110100010101011)) color_data = 12'b011111101110;
		if(({row_reg, col_reg}>=18'b010110100010101100) && ({row_reg, col_reg}<18'b010110100010111000)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010110100010111000) && ({row_reg, col_reg}<18'b010110100010111011)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010110100010111011)) color_data = 12'b101011101111;
		if(({row_reg, col_reg}==18'b010110100010111100)) color_data = 12'b101111101111;
		if(({row_reg, col_reg}==18'b010110100010111101)) color_data = 12'b011110011010;
		if(({row_reg, col_reg}==18'b010110100010111110)) color_data = 12'b010001110110;
		if(({row_reg, col_reg}==18'b010110100010111111)) color_data = 12'b010101110110;
		if(({row_reg, col_reg}==18'b010110100011000000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010110100011000001)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010110100011000010) && ({row_reg, col_reg}<18'b010110100011000101)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}>=18'b010110100011000101) && ({row_reg, col_reg}<18'b010110100011000111)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==18'b010110100011000111)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010110100011001000) && ({row_reg, col_reg}<18'b010110100011001100)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}==18'b010110100011001100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010110100011001101)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}>=18'b010110100011001110) && ({row_reg, col_reg}<18'b010110100011010000)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==18'b010110100011010000)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}>=18'b010110100011010001) && ({row_reg, col_reg}<18'b010110100011010011)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010110100011010011) && ({row_reg, col_reg}<18'b010110100011011010)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}>=18'b010110100011011010) && ({row_reg, col_reg}<18'b010110100011011110)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==18'b010110100011011110)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010110100011011111)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==18'b010110100011100000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010110100011100001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010110100011100010)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010110100011100011)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}>=18'b010110100011100100) && ({row_reg, col_reg}<18'b010110100011101001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010110100011101001)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}==18'b010110100011101010)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==18'b010110100011101011)) color_data = 12'b010101110111;
		if(({row_reg, col_reg}==18'b010110100011101100)) color_data = 12'b010101111001;
		if(({row_reg, col_reg}==18'b010110100011101101)) color_data = 12'b010001111001;
		if(({row_reg, col_reg}==18'b010110100011101110)) color_data = 12'b001101111010;
		if(({row_reg, col_reg}==18'b010110100011101111)) color_data = 12'b001110001011;
		if(({row_reg, col_reg}==18'b010110100011110000)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b010110100011110001)) color_data = 12'b010010101100;
		if(({row_reg, col_reg}==18'b010110100011110010)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010110100011110011) && ({row_reg, col_reg}<18'b010110100011110101)) color_data = 12'b100111111110;
		if(({row_reg, col_reg}==18'b010110100011110101)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010110100011110110) && ({row_reg, col_reg}<18'b010110100011111010)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010110100011111010)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010110100011111011)) color_data = 12'b010010101110;
		if(({row_reg, col_reg}>=18'b010110100011111100) && ({row_reg, col_reg}<18'b010110100011111110)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010110100011111110)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010110100011111111)) color_data = 12'b001110001011;
		if(({row_reg, col_reg}==18'b010110100100000000)) color_data = 12'b011111101111;
		if(({row_reg, col_reg}>=18'b010110100100000001) && ({row_reg, col_reg}<18'b010110100100000011)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}>=18'b010110100100000011) && ({row_reg, col_reg}<18'b010110100100000110)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010110100100000110)) color_data = 12'b100011111110;
		if(({row_reg, col_reg}==18'b010110100100000111)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010110100100001000)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010110100100001001)) color_data = 12'b011011001110;
		if(({row_reg, col_reg}==18'b010110100100001010)) color_data = 12'b001001111010;
		if(({row_reg, col_reg}>=18'b010110100100001011) && ({row_reg, col_reg}<18'b010110100100001101)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010110100100001101)) color_data = 12'b010001111101;
		if(({row_reg, col_reg}==18'b010110100100001110)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==18'b010110100100001111)) color_data = 12'b011010101111;

		if(({row_reg, col_reg}>=18'b010110100100010000) && ({row_reg, col_reg}<18'b010110101000010000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010110101000010000)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b010110101000010001)) color_data = 12'b010110011111;
		if(({row_reg, col_reg}>=18'b010110101000010010) && ({row_reg, col_reg}<18'b010110101000010110)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010110101000010110)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b010110101000010111) && ({row_reg, col_reg}<18'b010110101000011001)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}>=18'b010110101000011001) && ({row_reg, col_reg}<18'b010110101000011011)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010110101000011011)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}>=18'b010110101000011100) && ({row_reg, col_reg}<18'b010110101000011111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010110101000011111)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b010110101000100000) && ({row_reg, col_reg}<18'b010110101000100011)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b010110101000100011)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010110101000100100)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b010110101000100101)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010110101000100110)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}>=18'b010110101000100111) && ({row_reg, col_reg}<18'b010110101000101100)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b010110101000101100) && ({row_reg, col_reg}<18'b010110101000110000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010110101000110000)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b010110101000110001) && ({row_reg, col_reg}<18'b010110101000110011)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}>=18'b010110101000110011) && ({row_reg, col_reg}<18'b010110101000110110)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b010110101000110110)) color_data = 12'b011110111111;
		if(({row_reg, col_reg}==18'b010110101000110111)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b010110101000111000)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b010110101000111001) && ({row_reg, col_reg}<18'b010110101000111011)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b010110101000111011)) color_data = 12'b000101111010;
		if(({row_reg, col_reg}==18'b010110101000111100)) color_data = 12'b010010101100;
		if(({row_reg, col_reg}==18'b010110101000111101)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010110101000111110) && ({row_reg, col_reg}<18'b010110101001000011)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010110101001000011)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010110101001000100)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010110101001000101)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010110101001000110)) color_data = 12'b010010101101;
		if(({row_reg, col_reg}==18'b010110101001000111)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b010110101001001000) && ({row_reg, col_reg}<18'b010110101001001010)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010110101001001010) && ({row_reg, col_reg}<18'b010110101001001100)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b010110101001001100) && ({row_reg, col_reg}<18'b010110101001010000)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b010110101001010000) && ({row_reg, col_reg}<18'b010110101001010010)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010110101001010010)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010110101001010011)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b010110101001010100)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}>=18'b010110101001010101) && ({row_reg, col_reg}<18'b010110101001010111)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}>=18'b010110101001010111) && ({row_reg, col_reg}<18'b010110101001011001)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010110101001011001)) color_data = 12'b010010101100;
		if(({row_reg, col_reg}==18'b010110101001011010)) color_data = 12'b000101111011;
		if(({row_reg, col_reg}>=18'b010110101001011011) && ({row_reg, col_reg}<18'b010110101001011101)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b010110101001011101)) color_data = 12'b010001111010;
		if(({row_reg, col_reg}==18'b010110101001011110)) color_data = 12'b100010101011;
		if(({row_reg, col_reg}==18'b010110101001011111)) color_data = 12'b100110101011;
		if(({row_reg, col_reg}==18'b010110101001100000)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}>=18'b010110101001100001) && ({row_reg, col_reg}<18'b010110101001100100)) color_data = 12'b101110101001;
		if(({row_reg, col_reg}==18'b010110101001100100)) color_data = 12'b101010101001;
		if(({row_reg, col_reg}==18'b010110101001100101)) color_data = 12'b101010101010;
		if(({row_reg, col_reg}==18'b010110101001100110)) color_data = 12'b100110011010;
		if(({row_reg, col_reg}==18'b010110101001100111)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010110101001101000)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}>=18'b010110101001101001) && ({row_reg, col_reg}<18'b010110101001101011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010110101001101011) && ({row_reg, col_reg}<18'b010110101001101101)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}>=18'b010110101001101101) && ({row_reg, col_reg}<18'b010110101001101111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010110101001101111) && ({row_reg, col_reg}<18'b010110101001110001)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==18'b010110101001110001)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010110101001110010)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010110101001110011) && ({row_reg, col_reg}<18'b010110101001110101)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}>=18'b010110101001110101) && ({row_reg, col_reg}<18'b010110101001110111)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010110101001110111) && ({row_reg, col_reg}<18'b010110101001111010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010110101001111010)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010110101001111011)) color_data = 12'b101110101011;
		if(({row_reg, col_reg}>=18'b010110101001111100) && ({row_reg, col_reg}<18'b010110101001111110)) color_data = 12'b101010111100;
		if(({row_reg, col_reg}==18'b010110101001111110)) color_data = 12'b100110111101;
		if(({row_reg, col_reg}==18'b010110101001111111)) color_data = 12'b101011011110;
		if(({row_reg, col_reg}>=18'b010110101010000000) && ({row_reg, col_reg}<18'b010110101010000010)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}==18'b010110101010000010)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010110101010000011) && ({row_reg, col_reg}<18'b010110101010001000)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010110101010001000) && ({row_reg, col_reg}<18'b010110101010001101)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010110101010001101)) color_data = 12'b011011001110;
		if(({row_reg, col_reg}==18'b010110101010001110)) color_data = 12'b001110011011;
		if(({row_reg, col_reg}==18'b010110101010001111)) color_data = 12'b000101111011;
		if(({row_reg, col_reg}==18'b010110101010010000)) color_data = 12'b000101111100;
		if(({row_reg, col_reg}>=18'b010110101010010001) && ({row_reg, col_reg}<18'b010110101010010011)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010110101010010011)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010110101010010100)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b010110101010010101)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010110101010010110)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010110101010010111) && ({row_reg, col_reg}<18'b010110101010011001)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010110101010011001)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010110101010011010)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010110101010011011)) color_data = 12'b001110011100;
		if(({row_reg, col_reg}==18'b010110101010011100)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}>=18'b010110101010011101) && ({row_reg, col_reg}<18'b010110101010101011)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010110101010101011) && ({row_reg, col_reg}<18'b010110101010110000)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010110101010110000) && ({row_reg, col_reg}<18'b010110101010111000)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010110101010111000)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010110101010111001)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010110101010111010)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010110101010111011) && ({row_reg, col_reg}<18'b010110101010111101)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}==18'b010110101010111101)) color_data = 12'b011010101011;
		if(({row_reg, col_reg}==18'b010110101010111110)) color_data = 12'b001101110111;
		if(({row_reg, col_reg}==18'b010110101010111111)) color_data = 12'b010001110110;
		if(({row_reg, col_reg}==18'b010110101011000000)) color_data = 12'b010101110101;
		if(({row_reg, col_reg}>=18'b010110101011000001) && ({row_reg, col_reg}<18'b010110101011000011)) color_data = 12'b010101100101;
		if(({row_reg, col_reg}>=18'b010110101011000011) && ({row_reg, col_reg}<18'b010110101011000101)) color_data = 12'b010101110110;
		if(({row_reg, col_reg}>=18'b010110101011000101) && ({row_reg, col_reg}<18'b010110101011001000)) color_data = 12'b010101110111;
		if(({row_reg, col_reg}>=18'b010110101011001000) && ({row_reg, col_reg}<18'b010110101011001011)) color_data = 12'b010101110110;
		if(({row_reg, col_reg}==18'b010110101011001011)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}>=18'b010110101011001100) && ({row_reg, col_reg}<18'b010110101011001110)) color_data = 12'b010101110111;
		if(({row_reg, col_reg}==18'b010110101011001110)) color_data = 12'b011001111000;
		if(({row_reg, col_reg}==18'b010110101011001111)) color_data = 12'b010101100111;
		if(({row_reg, col_reg}==18'b010110101011010000)) color_data = 12'b010101111000;
		if(({row_reg, col_reg}>=18'b010110101011010001) && ({row_reg, col_reg}<18'b010110101011010011)) color_data = 12'b011001111000;
		if(({row_reg, col_reg}>=18'b010110101011010011) && ({row_reg, col_reg}<18'b010110101011010101)) color_data = 12'b010101101000;
		if(({row_reg, col_reg}==18'b010110101011010101)) color_data = 12'b011001101000;
		if(({row_reg, col_reg}==18'b010110101011010110)) color_data = 12'b011001111000;
		if(({row_reg, col_reg}>=18'b010110101011010111) && ({row_reg, col_reg}<18'b010110101011011101)) color_data = 12'b011001101000;
		if(({row_reg, col_reg}==18'b010110101011011101)) color_data = 12'b010101100111;
		if(({row_reg, col_reg}>=18'b010110101011011110) && ({row_reg, col_reg}<18'b010110101011100000)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}==18'b010110101011100000)) color_data = 12'b010101100110;
		if(({row_reg, col_reg}==18'b010110101011100001)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010110101011100010)) color_data = 12'b010101100110;
		if(({row_reg, col_reg}==18'b010110101011100011)) color_data = 12'b010101100111;
		if(({row_reg, col_reg}==18'b010110101011100100)) color_data = 12'b010101110111;
		if(({row_reg, col_reg}==18'b010110101011100101)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}>=18'b010110101011100110) && ({row_reg, col_reg}<18'b010110101011101000)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}==18'b010110101011101000)) color_data = 12'b010101100110;
		if(({row_reg, col_reg}==18'b010110101011101001)) color_data = 12'b010101110110;
		if(({row_reg, col_reg}==18'b010110101011101010)) color_data = 12'b010101110111;
		if(({row_reg, col_reg}==18'b010110101011101011)) color_data = 12'b010001111000;
		if(({row_reg, col_reg}==18'b010110101011101100)) color_data = 12'b010001111001;
		if(({row_reg, col_reg}>=18'b010110101011101101) && ({row_reg, col_reg}<18'b010110101011101111)) color_data = 12'b001101111010;
		if(({row_reg, col_reg}>=18'b010110101011101111) && ({row_reg, col_reg}<18'b010110101011110001)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b010110101011110001)) color_data = 12'b010010101100;
		if(({row_reg, col_reg}>=18'b010110101011110010) && ({row_reg, col_reg}<18'b010110101011111011)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010110101011111011)) color_data = 12'b001110011100;
		if(({row_reg, col_reg}==18'b010110101011111100)) color_data = 12'b000101111011;
		if(({row_reg, col_reg}==18'b010110101011111101)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b010110101011111110)) color_data = 12'b000101111010;
		if(({row_reg, col_reg}==18'b010110101011111111)) color_data = 12'b001110001010;
		if(({row_reg, col_reg}==18'b010110101100000000)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}>=18'b010110101100000001) && ({row_reg, col_reg}<18'b010110101100000110)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010110101100000110)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010110101100000111) && ({row_reg, col_reg}<18'b010110101100001001)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010110101100001001)) color_data = 12'b011011001111;
		if(({row_reg, col_reg}==18'b010110101100001010)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}>=18'b010110101100001011) && ({row_reg, col_reg}<18'b010110101100001101)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010110101100001101)) color_data = 12'b010001111101;
		if(({row_reg, col_reg}==18'b010110101100001110)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==18'b010110101100001111)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b010110101100010000)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b010110101100010001) && ({row_reg, col_reg}<18'b010110110000000100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010110110000000100)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010110110000000101) && ({row_reg, col_reg}<18'b010110110000000111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010110110000000111)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010110110000001000) && ({row_reg, col_reg}<18'b010110110000010000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010110110000010000)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b010110110000010001)) color_data = 12'b010110011111;
		if(({row_reg, col_reg}>=18'b010110110000010010) && ({row_reg, col_reg}<18'b010110110000010101)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010110110000010101)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010110110000010110)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b010110110000010111) && ({row_reg, col_reg}<18'b010110110000011100)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}>=18'b010110110000011100) && ({row_reg, col_reg}<18'b010110110000100000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010110110000100000)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010110110000100001)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010110110000100010) && ({row_reg, col_reg}<18'b010110110000100100)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010110110000100100)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}>=18'b010110110000100101) && ({row_reg, col_reg}<18'b010110110000100111)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b010110110000100111) && ({row_reg, col_reg}<18'b010110110000101001)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b010110110000101001) && ({row_reg, col_reg}<18'b010110110000101011)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010110110000101011)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010110110000101100)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010110110000101101)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010110110000101110)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}==18'b010110110000101111)) color_data = 12'b010010001110;
		if(({row_reg, col_reg}>=18'b010110110000110000) && ({row_reg, col_reg}<18'b010110110000110011)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}>=18'b010110110000110011) && ({row_reg, col_reg}<18'b010110110000110101)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}>=18'b010110110000110101) && ({row_reg, col_reg}<18'b010110110000110111)) color_data = 12'b010010011101;
		if(({row_reg, col_reg}==18'b010110110000110111)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}>=18'b010110110000111000) && ({row_reg, col_reg}<18'b010110110000111010)) color_data = 12'b010110101110;
		if(({row_reg, col_reg}==18'b010110110000111010)) color_data = 12'b010110111101;
		if(({row_reg, col_reg}==18'b010110110000111011)) color_data = 12'b010110101101;
		if(({row_reg, col_reg}==18'b010110110000111100)) color_data = 12'b010110111101;
		if(({row_reg, col_reg}>=18'b010110110000111101) && ({row_reg, col_reg}<18'b010110110001000100)) color_data = 12'b011011001110;
		if(({row_reg, col_reg}==18'b010110110001000100)) color_data = 12'b011011001111;
		if(({row_reg, col_reg}==18'b010110110001000101)) color_data = 12'b011010111111;
		if(({row_reg, col_reg}==18'b010110110001000110)) color_data = 12'b010010011101;
		if(({row_reg, col_reg}==18'b010110110001000111)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010110110001001000)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010110110001001001)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010110110001001010)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b010110110001001011) && ({row_reg, col_reg}<18'b010110110001001110)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b010110110001001110) && ({row_reg, col_reg}<18'b010110110001010000)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010110110001010000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010110110001010001)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010110110001010010)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010110110001010011)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010110110001010100)) color_data = 12'b010010011101;
		if(({row_reg, col_reg}==18'b010110110001010101)) color_data = 12'b011011001111;
		if(({row_reg, col_reg}>=18'b010110110001010110) && ({row_reg, col_reg}<18'b010110110001011001)) color_data = 12'b011011001110;
		if(({row_reg, col_reg}==18'b010110110001011001)) color_data = 12'b010110111101;
		if(({row_reg, col_reg}==18'b010110110001011010)) color_data = 12'b010010111101;
		if(({row_reg, col_reg}==18'b010110110001011011)) color_data = 12'b010110111101;
		if(({row_reg, col_reg}==18'b010110110001011100)) color_data = 12'b010110101101;
		if(({row_reg, col_reg}==18'b010110110001011101)) color_data = 12'b011010011011;
		if(({row_reg, col_reg}==18'b010110110001011110)) color_data = 12'b011110011010;
		if(({row_reg, col_reg}==18'b010110110001011111)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}==18'b010110110001100000)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==18'b010110110001100001)) color_data = 12'b100110000111;
		if(({row_reg, col_reg}>=18'b010110110001100010) && ({row_reg, col_reg}<18'b010110110001100101)) color_data = 12'b100110011000;
		if(({row_reg, col_reg}==18'b010110110001100101)) color_data = 12'b100110011001;
		if(({row_reg, col_reg}==18'b010110110001100110)) color_data = 12'b100010011001;
		if(({row_reg, col_reg}==18'b010110110001100111)) color_data = 12'b100010001001;
		if(({row_reg, col_reg}==18'b010110110001101000)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}==18'b010110110001101001)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010110110001101010)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010110110001101011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010110110001101100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010110110001101101) && ({row_reg, col_reg}<18'b010110110001101111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010110110001101111) && ({row_reg, col_reg}<18'b010110110001110010)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010110110001110010) && ({row_reg, col_reg}<18'b010110110001110100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010110110001110100) && ({row_reg, col_reg}<18'b010110110001110110)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010110110001110110) && ({row_reg, col_reg}<18'b010110110001111001)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010110110001111001)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==18'b010110110001111010)) color_data = 12'b011101111001;
		if(({row_reg, col_reg}==18'b010110110001111011)) color_data = 12'b100010001010;
		if(({row_reg, col_reg}>=18'b010110110001111100) && ({row_reg, col_reg}<18'b010110110001111110)) color_data = 12'b011110011011;
		if(({row_reg, col_reg}==18'b010110110001111110)) color_data = 12'b011010011100;
		if(({row_reg, col_reg}==18'b010110110001111111)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b010110110010000000) && ({row_reg, col_reg}<18'b010110110010000010)) color_data = 12'b011111001111;
		if(({row_reg, col_reg}>=18'b010110110010000010) && ({row_reg, col_reg}<18'b010110110010000100)) color_data = 12'b011011001111;
		if(({row_reg, col_reg}>=18'b010110110010000100) && ({row_reg, col_reg}<18'b010110110010001000)) color_data = 12'b011011011111;
		if(({row_reg, col_reg}>=18'b010110110010001000) && ({row_reg, col_reg}<18'b010110110010001100)) color_data = 12'b011011001110;
		if(({row_reg, col_reg}==18'b010110110010001100)) color_data = 12'b010111001110;
		if(({row_reg, col_reg}==18'b010110110010001101)) color_data = 12'b010110111110;
		if(({row_reg, col_reg}>=18'b010110110010001110) && ({row_reg, col_reg}<18'b010110110010010000)) color_data = 12'b010010101101;
		if(({row_reg, col_reg}==18'b010110110010010000)) color_data = 12'b010110101101;
		if(({row_reg, col_reg}==18'b010110110010010001)) color_data = 12'b010110111110;
		if(({row_reg, col_reg}==18'b010110110010010010)) color_data = 12'b010010011101;
		if(({row_reg, col_reg}==18'b010110110010010011)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010110110010010100)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010110110010010101) && ({row_reg, col_reg}<18'b010110110010010111)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010110110010010111)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b010110110010011000)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010110110010011001)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010110110010011010)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b010110110010011011)) color_data = 12'b001110011011;
		if(({row_reg, col_reg}==18'b010110110010011100)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}>=18'b010110110010011101) && ({row_reg, col_reg}<18'b010110110010101010)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010110110010101010)) color_data = 12'b011011011110;
		if(({row_reg, col_reg}==18'b010110110010101011)) color_data = 12'b010111001110;
		if(({row_reg, col_reg}>=18'b010110110010101100) && ({row_reg, col_reg}<18'b010110110010101111)) color_data = 12'b011011001110;
		if(({row_reg, col_reg}>=18'b010110110010101111) && ({row_reg, col_reg}<18'b010110110010111000)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010110110010111000)) color_data = 12'b011111101111;
		if(({row_reg, col_reg}==18'b010110110010111001)) color_data = 12'b010111001101;
		if(({row_reg, col_reg}==18'b010110110010111010)) color_data = 12'b011011001110;
		if(({row_reg, col_reg}>=18'b010110110010111011) && ({row_reg, col_reg}<18'b010110110010111101)) color_data = 12'b011011001101;
		if(({row_reg, col_reg}==18'b010110110010111101)) color_data = 12'b011010111100;
		if(({row_reg, col_reg}==18'b010110110010111110)) color_data = 12'b010110101010;
		if(({row_reg, col_reg}==18'b010110110010111111)) color_data = 12'b011010101001;
		if(({row_reg, col_reg}>=18'b010110110011000000) && ({row_reg, col_reg}<18'b010110110011000100)) color_data = 12'b011110101001;
		if(({row_reg, col_reg}==18'b010110110011000100)) color_data = 12'b011010011001;
		if(({row_reg, col_reg}==18'b010110110011000101)) color_data = 12'b011010101001;
		if(({row_reg, col_reg}==18'b010110110011000110)) color_data = 12'b011010011010;
		if(({row_reg, col_reg}==18'b010110110011000111)) color_data = 12'b011010011001;
		if(({row_reg, col_reg}==18'b010110110011001000)) color_data = 12'b011110101001;
		if(({row_reg, col_reg}==18'b010110110011001001)) color_data = 12'b011110011001;
		if(({row_reg, col_reg}==18'b010110110011001010)) color_data = 12'b011110101001;
		if(({row_reg, col_reg}==18'b010110110011001011)) color_data = 12'b011010011001;
		if(({row_reg, col_reg}==18'b010110110011001100)) color_data = 12'b010101111000;
		if(({row_reg, col_reg}>=18'b010110110011001101) && ({row_reg, col_reg}<18'b010110110011001111)) color_data = 12'b010101111001;
		if(({row_reg, col_reg}>=18'b010110110011001111) && ({row_reg, col_reg}<18'b010110110011010010)) color_data = 12'b010001111001;
		if(({row_reg, col_reg}>=18'b010110110011010010) && ({row_reg, col_reg}<18'b010110110011011101)) color_data = 12'b010101111001;
		if(({row_reg, col_reg}==18'b010110110011011101)) color_data = 12'b010001101000;
		if(({row_reg, col_reg}==18'b010110110011011110)) color_data = 12'b011010001001;
		if(({row_reg, col_reg}==18'b010110110011011111)) color_data = 12'b011110101011;
		if(({row_reg, col_reg}==18'b010110110011100000)) color_data = 12'b100010101001;
		if(({row_reg, col_reg}==18'b010110110011100001)) color_data = 12'b100010101010;
		if(({row_reg, col_reg}>=18'b010110110011100010) && ({row_reg, col_reg}<18'b010110110011101010)) color_data = 12'b011110011001;
		if(({row_reg, col_reg}==18'b010110110011101010)) color_data = 12'b011010011001;
		if(({row_reg, col_reg}==18'b010110110011101011)) color_data = 12'b011010011010;
		if(({row_reg, col_reg}==18'b010110110011101100)) color_data = 12'b011010011011;
		if(({row_reg, col_reg}==18'b010110110011101101)) color_data = 12'b010110101100;
		if(({row_reg, col_reg}>=18'b010110110011101110) && ({row_reg, col_reg}<18'b010110110011110000)) color_data = 12'b010110101101;
		if(({row_reg, col_reg}==18'b010110110011110000)) color_data = 12'b010010111101;
		if(({row_reg, col_reg}==18'b010110110011110001)) color_data = 12'b010111001101;
		if(({row_reg, col_reg}>=18'b010110110011110010) && ({row_reg, col_reg}<18'b010110110011111011)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010110110011111011)) color_data = 12'b010111001101;
		if(({row_reg, col_reg}==18'b010110110011111100)) color_data = 12'b010010101101;
		if(({row_reg, col_reg}==18'b010110110011111101)) color_data = 12'b010110111110;
		if(({row_reg, col_reg}==18'b010110110011111110)) color_data = 12'b010010101100;
		if(({row_reg, col_reg}==18'b010110110011111111)) color_data = 12'b010110111100;
		if(({row_reg, col_reg}>=18'b010110110100000000) && ({row_reg, col_reg}<18'b010110110100000110)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}>=18'b010110110100000110) && ({row_reg, col_reg}<18'b010110110100001000)) color_data = 12'b011011001110;
		if(({row_reg, col_reg}==18'b010110110100001000)) color_data = 12'b011011001111;
		if(({row_reg, col_reg}==18'b010110110100001001)) color_data = 12'b010110111110;
		if(({row_reg, col_reg}==18'b010110110100001010)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}>=18'b010110110100001011) && ({row_reg, col_reg}<18'b010110110100001101)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}==18'b010110110100001101)) color_data = 12'b010110001101;
		if(({row_reg, col_reg}==18'b010110110100001110)) color_data = 12'b011010011110;
		if(({row_reg, col_reg}==18'b010110110100001111)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b010110110100010000)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b010110110100010001) && ({row_reg, col_reg}<18'b010110111000000100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010110111000000100)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010110111000000101) && ({row_reg, col_reg}<18'b010110111000010000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010110111000010000)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b010110111000010001)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}>=18'b010110111000010010) && ({row_reg, col_reg}<18'b010110111000010110)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010110111000010110)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010110111000010111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010110111000011000) && ({row_reg, col_reg}<18'b010110111000011110)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}>=18'b010110111000011110) && ({row_reg, col_reg}<18'b010110111000100000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010110111000100000)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010110111000100001)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010110111000100010)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b010110111000100011) && ({row_reg, col_reg}<18'b010110111000100110)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010110111000100110)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010110111000100111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010110111000101000) && ({row_reg, col_reg}<18'b010110111000101101)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010110111000101101)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b010110111000101110)) color_data = 12'b010010011110;
		if(({row_reg, col_reg}==18'b010110111000101111)) color_data = 12'b010110101111;
		if(({row_reg, col_reg}>=18'b010110111000110000) && ({row_reg, col_reg}<18'b010110111000110010)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b010110111000110010)) color_data = 12'b011010111111;
		if(({row_reg, col_reg}>=18'b010110111000110011) && ({row_reg, col_reg}<18'b010110111000110101)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010110111000110101)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010110111000110110)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010110111000110111)) color_data = 12'b010010011101;
		if(({row_reg, col_reg}==18'b010110111000111000)) color_data = 12'b100011011111;
		if(({row_reg, col_reg}==18'b010110111000111001)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b010110111000111010)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010110111000111011)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b010110111000111100)) color_data = 12'b011111001111;
		if(({row_reg, col_reg}==18'b010110111000111101)) color_data = 12'b001110011100;
		if(({row_reg, col_reg}>=18'b010110111000111110) && ({row_reg, col_reg}<18'b010110111001000010)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b010110111001000010)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b010110111001000011)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b010110111001000100)) color_data = 12'b001010001101;
		if(({row_reg, col_reg}==18'b010110111001000101)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}>=18'b010110111001000110) && ({row_reg, col_reg}<18'b010110111001001000)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010110111001001000)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}>=18'b010110111001001001) && ({row_reg, col_reg}<18'b010110111001001011)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010110111001001011) && ({row_reg, col_reg}<18'b010110111001001111)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010110111001001111)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}>=18'b010110111001010000) && ({row_reg, col_reg}<18'b010110111001010011)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010110111001010011)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010110111001010100)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b010110111001010101) && ({row_reg, col_reg}<18'b010110111001010111)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}>=18'b010110111001010111) && ({row_reg, col_reg}<18'b010110111001011001)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b010110111001011001)) color_data = 12'b011011001110;
		if(({row_reg, col_reg}>=18'b010110111001011010) && ({row_reg, col_reg}<18'b010110111001011100)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010110111001011100)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}==18'b010110111001011101)) color_data = 12'b100111011110;
		if(({row_reg, col_reg}==18'b010110111001011110)) color_data = 12'b011110101010;
		if(({row_reg, col_reg}==18'b010110111001011111)) color_data = 12'b011010000111;
		if(({row_reg, col_reg}==18'b010110111001100000)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010110111001100001)) color_data = 12'b011110000110;
		if(({row_reg, col_reg}==18'b010110111001100010)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010110111001100011)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010110111001100100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010110111001100101)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==18'b010110111001100110)) color_data = 12'b100010001000;
		if(({row_reg, col_reg}==18'b010110111001100111)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==18'b010110111001101000)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010110111001101001)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010110111001101010)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010110111001101011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010110111001101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010110111001101101) && ({row_reg, col_reg}<18'b010110111001101111)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}>=18'b010110111001101111) && ({row_reg, col_reg}<18'b010110111001110010)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==18'b010110111001110010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010110111001110011) && ({row_reg, col_reg}<18'b010110111001111000)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010110111001111000)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010110111001111001)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}==18'b010110111001111010)) color_data = 12'b011001111001;
		if(({row_reg, col_reg}==18'b010110111001111011)) color_data = 12'b011001111010;
		if(({row_reg, col_reg}==18'b010110111001111100)) color_data = 12'b010101111011;
		if(({row_reg, col_reg}==18'b010110111001111101)) color_data = 12'b010001111011;
		if(({row_reg, col_reg}>=18'b010110111001111110) && ({row_reg, col_reg}<18'b010110111010000000)) color_data = 12'b001101111011;
		if(({row_reg, col_reg}>=18'b010110111010000000) && ({row_reg, col_reg}<18'b010110111010000010)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b010110111010000010)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b010110111010000011)) color_data = 12'b000110001100;
		if(({row_reg, col_reg}==18'b010110111010000100)) color_data = 12'b000101111100;
		if(({row_reg, col_reg}==18'b010110111010000101)) color_data = 12'b000110001100;
		if(({row_reg, col_reg}==18'b010110111010000110)) color_data = 12'b000101111100;
		if(({row_reg, col_reg}==18'b010110111010000111)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b010110111010001000) && ({row_reg, col_reg}<18'b010110111010001100)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b010110111010001100)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b010110111010001101)) color_data = 12'b010010101101;
		if(({row_reg, col_reg}==18'b010110111010001110)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}>=18'b010110111010001111) && ({row_reg, col_reg}<18'b010110111010010001)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010110111010010001)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010110111010010010)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==18'b010110111010010011)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010110111010010100)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010110111010010101)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b010110111010010110) && ({row_reg, col_reg}<18'b010110111010011000)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b010110111010011000)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010110111010011001)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010110111010011010)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b010110111010011011)) color_data = 12'b001110011011;
		if(({row_reg, col_reg}==18'b010110111010011100)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}>=18'b010110111010011101) && ({row_reg, col_reg}<18'b010110111010100110)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010110111010100110)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010110111010100111) && ({row_reg, col_reg}<18'b010110111010101001)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010110111010101001)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010110111010101010)) color_data = 12'b010110111101;
		if(({row_reg, col_reg}>=18'b010110111010101011) && ({row_reg, col_reg}<18'b010110111010101101)) color_data = 12'b000101111011;
		if(({row_reg, col_reg}==18'b010110111010101101)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b010110111010101110)) color_data = 12'b001110011011;
		if(({row_reg, col_reg}==18'b010110111010101111)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}>=18'b010110111010110000) && ({row_reg, col_reg}<18'b010110111010111000)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010110111010111000)) color_data = 12'b011011001101;
		if(({row_reg, col_reg}==18'b010110111010111001)) color_data = 12'b001010001010;
		if(({row_reg, col_reg}==18'b010110111010111010)) color_data = 12'b001010011011;
		if(({row_reg, col_reg}==18'b010110111010111011)) color_data = 12'b001010001010;
		if(({row_reg, col_reg}==18'b010110111010111100)) color_data = 12'b001110011010;
		if(({row_reg, col_reg}==18'b010110111010111101)) color_data = 12'b011010111100;
		if(({row_reg, col_reg}==18'b010110111010111110)) color_data = 12'b100111101110;
		if(({row_reg, col_reg}==18'b010110111010111111)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}==18'b010110111011000000)) color_data = 12'b101111101110;
		if(({row_reg, col_reg}>=18'b010110111011000001) && ({row_reg, col_reg}<18'b010110111011000011)) color_data = 12'b101011101110;
		if(({row_reg, col_reg}==18'b010110111011000011)) color_data = 12'b101111111110;
		if(({row_reg, col_reg}>=18'b010110111011000100) && ({row_reg, col_reg}<18'b010110111011001001)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}==18'b010110111011001001)) color_data = 12'b101111111111;
		if(({row_reg, col_reg}==18'b010110111011001010)) color_data = 12'b101111101111;
		if(({row_reg, col_reg}==18'b010110111011001011)) color_data = 12'b011110111100;
		if(({row_reg, col_reg}>=18'b010110111011001100) && ({row_reg, col_reg}<18'b010110111011001111)) color_data = 12'b010001111010;
		if(({row_reg, col_reg}==18'b010110111011001111)) color_data = 12'b001101111010;
		if(({row_reg, col_reg}>=18'b010110111011010000) && ({row_reg, col_reg}<18'b010110111011011010)) color_data = 12'b010001111011;
		if(({row_reg, col_reg}>=18'b010110111011011010) && ({row_reg, col_reg}<18'b010110111011011101)) color_data = 12'b010001111010;
		if(({row_reg, col_reg}==18'b010110111011011101)) color_data = 12'b001101111001;
		if(({row_reg, col_reg}==18'b010110111011011110)) color_data = 12'b011010101100;
		if(({row_reg, col_reg}==18'b010110111011011111)) color_data = 12'b100111011111;
		if(({row_reg, col_reg}>=18'b010110111011100000) && ({row_reg, col_reg}<18'b010110111011100011)) color_data = 12'b101011101110;
		if(({row_reg, col_reg}>=18'b010110111011100011) && ({row_reg, col_reg}<18'b010110111011101000)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}==18'b010110111011101000)) color_data = 12'b101011111110;
		if(({row_reg, col_reg}>=18'b010110111011101001) && ({row_reg, col_reg}<18'b010110111011101101)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}>=18'b010110111011101101) && ({row_reg, col_reg}<18'b010110111011110000)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010110111011110000) && ({row_reg, col_reg}<18'b010110111011111101)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010110111011111101) && ({row_reg, col_reg}<18'b010110111011111111)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010110111011111111)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010110111100000000)) color_data = 12'b011111001110;
		if(({row_reg, col_reg}==18'b010110111100000001)) color_data = 12'b010110111101;
		if(({row_reg, col_reg}>=18'b010110111100000010) && ({row_reg, col_reg}<18'b010110111100000100)) color_data = 12'b010110111110;
		if(({row_reg, col_reg}==18'b010110111100000100)) color_data = 12'b010010011101;
		if(({row_reg, col_reg}==18'b010110111100000101)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}>=18'b010110111100000110) && ({row_reg, col_reg}<18'b010110111100001000)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b010110111100001000)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b010110111100001001)) color_data = 12'b010010011101;
		if(({row_reg, col_reg}==18'b010110111100001010)) color_data = 12'b010110101110;
		if(({row_reg, col_reg}>=18'b010110111100001011) && ({row_reg, col_reg}<18'b010110111100010000)) color_data = 12'b011010101111;

		if(({row_reg, col_reg}>=18'b010110111100010000) && ({row_reg, col_reg}<18'b010111000000010000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010111000000010000)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b010111000000010001)) color_data = 12'b011010011110;
		if(({row_reg, col_reg}>=18'b010111000000010010) && ({row_reg, col_reg}<18'b010111000000010100)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}>=18'b010111000000010100) && ({row_reg, col_reg}<18'b010111000000010111)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010111000000010111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010111000000011000) && ({row_reg, col_reg}<18'b010111000000011101)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}>=18'b010111000000011101) && ({row_reg, col_reg}<18'b010111000000100101)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111000000100101)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b010111000000100110) && ({row_reg, col_reg}<18'b010111000000101001)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010111000000101001) && ({row_reg, col_reg}<18'b010111000000101011)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b010111000000101011) && ({row_reg, col_reg}<18'b010111000000101101)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111000000101101)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010111000000101110)) color_data = 12'b010010011110;
		if(({row_reg, col_reg}>=18'b010111000000101111) && ({row_reg, col_reg}<18'b010111000000110010)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b010111000000110010)) color_data = 12'b010110101111;
		if(({row_reg, col_reg}==18'b010111000000110011)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}==18'b010111000000110100)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b010111000000110101)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010111000000110110)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b010111000000110111)) color_data = 12'b010010011100;
		if(({row_reg, col_reg}==18'b010111000000111000)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010111000000111001)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}==18'b010111000000111010)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b010111000000111011)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010111000000111100)) color_data = 12'b011111001111;
		if(({row_reg, col_reg}==18'b010111000000111101)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b010111000000111110)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}>=18'b010111000000111111) && ({row_reg, col_reg}<18'b010111000001000001)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b010111000001000001)) color_data = 12'b001010001101;
		if(({row_reg, col_reg}>=18'b010111000001000010) && ({row_reg, col_reg}<18'b010111000001001000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010111000001001000) && ({row_reg, col_reg}<18'b010111000001001010)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010111000001001010)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111000001001011)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b010111000001001100) && ({row_reg, col_reg}<18'b010111000001001110)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b010111000001001110)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010111000001001111)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b010111000001010000)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b010111000001010001) && ({row_reg, col_reg}<18'b010111000001010011)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010111000001010011)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b010111000001010100) && ({row_reg, col_reg}<18'b010111000001010110)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111000001010110)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b010111000001010111)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b010111000001011000)) color_data = 12'b000101111011;
		if(({row_reg, col_reg}==18'b010111000001011001)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}==18'b010111000001011010)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010111000001011011)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010111000001011100)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}==18'b010111000001011101)) color_data = 12'b101011101110;
		if(({row_reg, col_reg}==18'b010111000001011110)) color_data = 12'b011010011001;
		if(({row_reg, col_reg}==18'b010111000001011111)) color_data = 12'b010101110111;
		if(({row_reg, col_reg}==18'b010111000001100000)) color_data = 12'b011110000111;
		if(({row_reg, col_reg}==18'b010111000001100001)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010111000001100010)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010111000001100011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010111000001100100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010111000001100101) && ({row_reg, col_reg}<18'b010111000001100111)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}==18'b010111000001100111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010111000001101000)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010111000001101001) && ({row_reg, col_reg}<18'b010111000001101101)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010111000001101101)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}>=18'b010111000001101110) && ({row_reg, col_reg}<18'b010111000001110011)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010111000001110011)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}==18'b010111000001110100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010111000001110101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010111000001110110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010111000001110111)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010111000001111000)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}==18'b010111000001111001)) color_data = 12'b010101101000;
		if(({row_reg, col_reg}==18'b010111000001111010)) color_data = 12'b010101111010;
		if(({row_reg, col_reg}==18'b010111000001111011)) color_data = 12'b010101111011;
		if(({row_reg, col_reg}==18'b010111000001111100)) color_data = 12'b010001111100;
		if(({row_reg, col_reg}>=18'b010111000001111101) && ({row_reg, col_reg}<18'b010111000001111111)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010111000001111111)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b010111000010000000) && ({row_reg, col_reg}<18'b010111000010000100)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010111000010000100) && ({row_reg, col_reg}<18'b010111000010000110)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b010111000010000110)) color_data = 12'b001010001110;
		if(({row_reg, col_reg}==18'b010111000010000111)) color_data = 12'b001010001101;
		if(({row_reg, col_reg}==18'b010111000010001000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010111000010001001) && ({row_reg, col_reg}<18'b010111000010001011)) color_data = 12'b001010001101;
		if(({row_reg, col_reg}==18'b010111000010001011)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111000010001100)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b010111000010001101)) color_data = 12'b010010101101;
		if(({row_reg, col_reg}>=18'b010111000010001110) && ({row_reg, col_reg}<18'b010111000010010010)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010111000010010010)) color_data = 12'b010110101101;
		if(({row_reg, col_reg}==18'b010111000010010011)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b010111000010010100) && ({row_reg, col_reg}<18'b010111000010011000)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b010111000010011000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111000010011001)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b010111000010011010)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b010111000010011011)) color_data = 12'b001110011011;
		if(({row_reg, col_reg}==18'b010111000010011100)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}>=18'b010111000010011101) && ({row_reg, col_reg}<18'b010111000010100101)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010111000010100101)) color_data = 12'b100011101110;
		if(({row_reg, col_reg}==18'b010111000010100110)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010111000010100111) && ({row_reg, col_reg}<18'b010111000010101001)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010111000010101001)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010111000010101010)) color_data = 12'b010010101100;
		if(({row_reg, col_reg}>=18'b010111000010101011) && ({row_reg, col_reg}<18'b010111000010101111)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b010111000010101111)) color_data = 12'b011111101111;
		if(({row_reg, col_reg}>=18'b010111000010110000) && ({row_reg, col_reg}<18'b010111000010110010)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010111000010110010)) color_data = 12'b011111111111;
		if(({row_reg, col_reg}>=18'b010111000010110011) && ({row_reg, col_reg}<18'b010111000010110111)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010111000010110111)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010111000010111000)) color_data = 12'b010110111101;
		if(({row_reg, col_reg}>=18'b010111000010111001) && ({row_reg, col_reg}<18'b010111000010111011)) color_data = 12'b000101111010;
		if(({row_reg, col_reg}>=18'b010111000010111011) && ({row_reg, col_reg}<18'b010111000010111101)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b010111000010111101)) color_data = 12'b011011001110;
		if(({row_reg, col_reg}>=18'b010111000010111110) && ({row_reg, col_reg}<18'b010111000011000011)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}>=18'b010111000011000011) && ({row_reg, col_reg}<18'b010111000011001000)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010111000011001000)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b010111000011001001)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}==18'b010111000011001010)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b010111000011001011)) color_data = 12'b011111001110;
		if(({row_reg, col_reg}>=18'b010111000011001100) && ({row_reg, col_reg}<18'b010111000011010000)) color_data = 12'b001101111011;
		if(({row_reg, col_reg}==18'b010111000011010000)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}>=18'b010111000011010001) && ({row_reg, col_reg}<18'b010111000011010011)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010111000011010011)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b010111000011010100) && ({row_reg, col_reg}<18'b010111000011010110)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010111000011010110)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b010111000011010111) && ({row_reg, col_reg}<18'b010111000011011011)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}>=18'b010111000011011011) && ({row_reg, col_reg}<18'b010111000011011101)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b010111000011011101)) color_data = 12'b001001111010;
		if(({row_reg, col_reg}==18'b010111000011011110)) color_data = 12'b010010101101;
		if(({row_reg, col_reg}==18'b010111000011011111)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}>=18'b010111000011100000) && ({row_reg, col_reg}<18'b010111000011100010)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010111000011100010) && ({row_reg, col_reg}<18'b010111000011100111)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010111000011100111) && ({row_reg, col_reg}<18'b010111000011101100)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010111000011101100) && ({row_reg, col_reg}<18'b010111000011110010)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010111000011110010)) color_data = 12'b011111111111;
		if(({row_reg, col_reg}>=18'b010111000011110011) && ({row_reg, col_reg}<18'b010111000011111001)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010111000011111001) && ({row_reg, col_reg}<18'b010111000011111101)) color_data = 12'b100011111110;
		if(({row_reg, col_reg}>=18'b010111000011111101) && ({row_reg, col_reg}<18'b010111000011111111)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010111000011111111)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010111000100000000) && ({row_reg, col_reg}<18'b010111000100000010)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==18'b010111000100000010)) color_data = 12'b011010111111;
		if(({row_reg, col_reg}==18'b010111000100000011)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b010111000100000100)) color_data = 12'b010010011110;
		if(({row_reg, col_reg}==18'b010111000100000101)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}>=18'b010111000100000110) && ({row_reg, col_reg}<18'b010111000100001000)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010111000100001000)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b010111000100001001)) color_data = 12'b001110011101;
		if(({row_reg, col_reg}==18'b010111000100001010)) color_data = 12'b011010111111;
		if(({row_reg, col_reg}==18'b010111000100001011)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b010111000100001100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010111000100001101)) color_data = 12'b011110101111;

		if(({row_reg, col_reg}>=18'b010111000100001110) && ({row_reg, col_reg}<18'b010111001000010000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010111001000010000)) color_data = 12'b011110111111;
		if(({row_reg, col_reg}==18'b010111001000010001)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==18'b010111001000010010)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}>=18'b010111001000010011) && ({row_reg, col_reg}<18'b010111001000010101)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b010111001000010101) && ({row_reg, col_reg}<18'b010111001000010111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111001000010111)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010111001000011000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111001000011001)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010111001000011010)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111001000011011)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b010111001000011100)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010111001000011101)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111001000011110)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010111001000011111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010111001000100000) && ({row_reg, col_reg}<18'b010111001000100100)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b010111001000100100) && ({row_reg, col_reg}<18'b010111001000101000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111001000101000)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010111001000101001)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111001000101010)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010111001000101011)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010111001000101100)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010111001000101101)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b010111001000101110)) color_data = 12'b010010011110;
		if(({row_reg, col_reg}>=18'b010111001000101111) && ({row_reg, col_reg}<18'b010111001000110010)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b010111001000110010)) color_data = 12'b010110101111;
		if(({row_reg, col_reg}==18'b010111001000110011)) color_data = 12'b010010001110;
		if(({row_reg, col_reg}==18'b010111001000110100)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010111001000110101)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111001000110110)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010111001000110111)) color_data = 12'b001110011100;
		if(({row_reg, col_reg}==18'b010111001000111000)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b010111001000111001)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010111001000111010) && ({row_reg, col_reg}<18'b010111001000111100)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b010111001000111100)) color_data = 12'b011011001111;
		if(({row_reg, col_reg}==18'b010111001000111101)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}>=18'b010111001000111110) && ({row_reg, col_reg}<18'b010111001001000000)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b010111001001000000)) color_data = 12'b001010001101;
		if(({row_reg, col_reg}==18'b010111001001000001)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010111001001000010)) color_data = 12'b000101111100;
		if(({row_reg, col_reg}>=18'b010111001001000011) && ({row_reg, col_reg}<18'b010111001001000101)) color_data = 12'b001010001101;
		if(({row_reg, col_reg}>=18'b010111001001000101) && ({row_reg, col_reg}<18'b010111001001000111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111001001000111)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b010111001001001000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111001001001001)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}>=18'b010111001001001010) && ({row_reg, col_reg}<18'b010111001001001101)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010111001001001101) && ({row_reg, col_reg}<18'b010111001001010000)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}>=18'b010111001001010000) && ({row_reg, col_reg}<18'b010111001001010010)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b010111001001010010)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b010111001001010011) && ({row_reg, col_reg}<18'b010111001001010101)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}>=18'b010111001001010101) && ({row_reg, col_reg}<18'b010111001001010111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111001001010111)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010111001001011000)) color_data = 12'b000101111010;
		if(({row_reg, col_reg}==18'b010111001001011001)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}==18'b010111001001011010)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010111001001011011) && ({row_reg, col_reg}<18'b010111001001011101)) color_data = 12'b100111111110;
		if(({row_reg, col_reg}==18'b010111001001011101)) color_data = 12'b101011101110;
		if(({row_reg, col_reg}==18'b010111001001011110)) color_data = 12'b010110011001;
		if(({row_reg, col_reg}==18'b010111001001011111)) color_data = 12'b010110001000;
		if(({row_reg, col_reg}>=18'b010111001001100000) && ({row_reg, col_reg}<18'b010111001001100010)) color_data = 12'b011110001000;
		if(({row_reg, col_reg}==18'b010111001001100010)) color_data = 12'b011101111000;
		if(({row_reg, col_reg}>=18'b010111001001100011) && ({row_reg, col_reg}<18'b010111001001100110)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}==18'b010111001001100110)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}>=18'b010111001001100111) && ({row_reg, col_reg}<18'b010111001001101011)) color_data = 12'b100010000111;
		if(({row_reg, col_reg}==18'b010111001001101011)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010111001001101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010111001001101101) && ({row_reg, col_reg}<18'b010111001001110010)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010111001001110010) && ({row_reg, col_reg}<18'b010111001001110100)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}>=18'b010111001001110100) && ({row_reg, col_reg}<18'b010111001001110110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010111001001110110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010111001001110111)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==18'b010111001001111000)) color_data = 12'b011001111000;
		if(({row_reg, col_reg}==18'b010111001001111001)) color_data = 12'b010001101001;
		if(({row_reg, col_reg}==18'b010111001001111010)) color_data = 12'b010001111010;
		if(({row_reg, col_reg}==18'b010111001001111011)) color_data = 12'b010001111011;
		if(({row_reg, col_reg}==18'b010111001001111100)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}>=18'b010111001001111101) && ({row_reg, col_reg}<18'b010111001010000000)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b010111001010000000) && ({row_reg, col_reg}<18'b010111001010000011)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b010111001010000011) && ({row_reg, col_reg}<18'b010111001010000111)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b010111001010000111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111001010001000)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}>=18'b010111001010001001) && ({row_reg, col_reg}<18'b010111001010001011)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111001010001011)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}==18'b010111001010001100)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b010111001010001101)) color_data = 12'b010010011101;
		if(({row_reg, col_reg}==18'b010111001010001110)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b010111001010001111)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}>=18'b010111001010010000) && ({row_reg, col_reg}<18'b010111001010010010)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010111001010010010)) color_data = 12'b010110111110;
		if(({row_reg, col_reg}==18'b010111001010010011)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010111001010010100)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b010111001010010101)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b010111001010010110) && ({row_reg, col_reg}<18'b010111001010011000)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b010111001010011000)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010111001010011001)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111001010011010)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b010111001010011011)) color_data = 12'b001110011100;
		if(({row_reg, col_reg}==18'b010111001010011100)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}>=18'b010111001010011101) && ({row_reg, col_reg}<18'b010111001010100001)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010111001010100001)) color_data = 12'b100011111110;
		if(({row_reg, col_reg}==18'b010111001010100010)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010111001010100011)) color_data = 12'b100011111110;
		if(({row_reg, col_reg}==18'b010111001010100100)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010111001010100101)) color_data = 12'b100011111110;
		if(({row_reg, col_reg}==18'b010111001010100110)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010111001010100111) && ({row_reg, col_reg}<18'b010111001010101001)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010111001010101001)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010111001010101010)) color_data = 12'b010010101100;
		if(({row_reg, col_reg}==18'b010111001010101011)) color_data = 12'b001010001010;
		if(({row_reg, col_reg}>=18'b010111001010101100) && ({row_reg, col_reg}<18'b010111001010101111)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b010111001010101111)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}>=18'b010111001010110000) && ({row_reg, col_reg}<18'b010111001010110110)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010111001010110110) && ({row_reg, col_reg}<18'b010111001010111000)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010111001010111000)) color_data = 12'b011111001111;
		if(({row_reg, col_reg}==18'b010111001010111001)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}>=18'b010111001010111010) && ({row_reg, col_reg}<18'b010111001010111100)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b010111001010111100)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b010111001010111101)) color_data = 12'b011011001110;
		if(({row_reg, col_reg}==18'b010111001010111110)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010111001010111111)) color_data = 12'b100011101110;
		if(({row_reg, col_reg}>=18'b010111001011000000) && ({row_reg, col_reg}<18'b010111001011000101)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010111001011000101) && ({row_reg, col_reg}<18'b010111001011001000)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010111001011001000) && ({row_reg, col_reg}<18'b010111001011001011)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010111001011001011)) color_data = 12'b011111001111;
		if(({row_reg, col_reg}==18'b010111001011001100)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b010111001011001101)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010111001011001110)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b010111001011001111)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010111001011010000)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}>=18'b010111001011010001) && ({row_reg, col_reg}<18'b010111001011011000)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010111001011011000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111001011011001)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010111001011011010)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010111001011011011) && ({row_reg, col_reg}<18'b010111001011011101)) color_data = 12'b001010001101;
		if(({row_reg, col_reg}==18'b010111001011011101)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b010111001011011110)) color_data = 12'b010010111110;
		if(({row_reg, col_reg}>=18'b010111001011011111) && ({row_reg, col_reg}<18'b010111001011111001)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010111001011111001) && ({row_reg, col_reg}<18'b010111001011111100)) color_data = 12'b100011111110;
		if(({row_reg, col_reg}>=18'b010111001011111100) && ({row_reg, col_reg}<18'b010111001011111110)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010111001011111110) && ({row_reg, col_reg}<18'b010111001100000000)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}>=18'b010111001100000000) && ({row_reg, col_reg}<18'b010111001100000010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010111001100000010) && ({row_reg, col_reg}<18'b010111001100000100)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b010111001100000100)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==18'b010111001100000101)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}>=18'b010111001100000110) && ({row_reg, col_reg}<18'b010111001100001000)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b010111001100001000)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010111001100001001)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}>=18'b010111001100001010) && ({row_reg, col_reg}<18'b010111001100010010)) color_data = 12'b011010101110;

		if(({row_reg, col_reg}==18'b010111001100010010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010111010000000000) && ({row_reg, col_reg}<18'b010111010000010000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010111010000010000)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}==18'b010111010000010001)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==18'b010111010000010010)) color_data = 12'b010001111100;
		if(({row_reg, col_reg}==18'b010111010000010011)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}>=18'b010111010000010100) && ({row_reg, col_reg}<18'b010111010000011001)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b010111010000011001) && ({row_reg, col_reg}<18'b010111010000011100)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010111010000011100)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010111010000011101)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111010000011110)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b010111010000011111) && ({row_reg, col_reg}<18'b010111010000100100)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111010000100100)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}>=18'b010111010000100101) && ({row_reg, col_reg}<18'b010111010000101010)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010111010000101010) && ({row_reg, col_reg}<18'b010111010000101100)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b010111010000101100)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111010000101101)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010111010000101110)) color_data = 12'b010010011110;
		if(({row_reg, col_reg}>=18'b010111010000101111) && ({row_reg, col_reg}<18'b010111010000110011)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b010111010000110011)) color_data = 12'b010010001110;
		if(({row_reg, col_reg}>=18'b010111010000110100) && ({row_reg, col_reg}<18'b010111010000110110)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111010000110110)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010111010000110111)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b010111010000111000)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010111010000111001)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010111010000111010)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b010111010000111011)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010111010000111100)) color_data = 12'b011011001111;
		if(({row_reg, col_reg}==18'b010111010000111101)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b010111010000111110)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}>=18'b010111010000111111) && ({row_reg, col_reg}<18'b010111010001000001)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}>=18'b010111010001000001) && ({row_reg, col_reg}<18'b010111010001001000)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b010111010001001000)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}>=18'b010111010001001001) && ({row_reg, col_reg}<18'b010111010001010000)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}>=18'b010111010001010000) && ({row_reg, col_reg}<18'b010111010001010100)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}>=18'b010111010001010100) && ({row_reg, col_reg}<18'b010111010001010110)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b010111010001010110)) color_data = 12'b001010001101;
		if(({row_reg, col_reg}==18'b010111010001010111)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b010111010001011000)) color_data = 12'b001010001010;
		if(({row_reg, col_reg}==18'b010111010001011001)) color_data = 12'b011111101111;
		if(({row_reg, col_reg}>=18'b010111010001011010) && ({row_reg, col_reg}<18'b010111010001011101)) color_data = 12'b100011111110;
		if(({row_reg, col_reg}==18'b010111010001011101)) color_data = 12'b100111101110;
		if(({row_reg, col_reg}==18'b010111010001011110)) color_data = 12'b011010101010;
		if(({row_reg, col_reg}==18'b010111010001011111)) color_data = 12'b010110001010;
		if(({row_reg, col_reg}>=18'b010111010001100000) && ({row_reg, col_reg}<18'b010111010001100010)) color_data = 12'b011110001010;
		if(({row_reg, col_reg}==18'b010111010001100010)) color_data = 12'b100001111001;
		if(({row_reg, col_reg}==18'b010111010001100011)) color_data = 12'b100001111000;
		if(({row_reg, col_reg}>=18'b010111010001100100) && ({row_reg, col_reg}<18'b010111010001101000)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010111010001101000)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}>=18'b010111010001101001) && ({row_reg, col_reg}<18'b010111010001101100)) color_data = 12'b100001110111;
		if(({row_reg, col_reg}==18'b010111010001101100)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}>=18'b010111010001101101) && ({row_reg, col_reg}<18'b010111010001101111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010111010001101111) && ({row_reg, col_reg}<18'b010111010001110010)) color_data = 12'b100001100110;
		if(({row_reg, col_reg}>=18'b010111010001110010) && ({row_reg, col_reg}<18'b010111010001110100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010111010001110100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}==18'b010111010001110101)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==18'b010111010001110110)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}==18'b010111010001110111)) color_data = 12'b011001111000;
		if(({row_reg, col_reg}==18'b010111010001111000)) color_data = 12'b010101111001;
		if(({row_reg, col_reg}==18'b010111010001111001)) color_data = 12'b010001111001;
		if(({row_reg, col_reg}==18'b010111010001111010)) color_data = 12'b010010001011;
		if(({row_reg, col_reg}>=18'b010111010001111011) && ({row_reg, col_reg}<18'b010111010001111101)) color_data = 12'b001110001011;
		if(({row_reg, col_reg}==18'b010111010001111101)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}>=18'b010111010001111110) && ({row_reg, col_reg}<18'b010111010010000000)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b010111010010000000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010111010010000001) && ({row_reg, col_reg}<18'b010111010010000110)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b010111010010000110) && ({row_reg, col_reg}<18'b010111010010001000)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010111010010001000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111010010001001)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}>=18'b010111010010001010) && ({row_reg, col_reg}<18'b010111010010001101)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111010010001101)) color_data = 12'b010010101110;
		if(({row_reg, col_reg}==18'b010111010010001110)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010111010010001111)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b010111010010010000)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010111010010010001)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b010111010010010010)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}>=18'b010111010010010011) && ({row_reg, col_reg}<18'b010111010010010101)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010111010010010101) && ({row_reg, col_reg}<18'b010111010010011000)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}>=18'b010111010010011000) && ({row_reg, col_reg}<18'b010111010010011010)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111010010011010)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010111010010011011)) color_data = 12'b001110011101;
		if(({row_reg, col_reg}==18'b010111010010011100)) color_data = 12'b100011011111;
		if(({row_reg, col_reg}==18'b010111010010011101)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010111010010011110)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010111010010011111)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}>=18'b010111010010100000) && ({row_reg, col_reg}<18'b010111010010100111)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010111010010100111)) color_data = 12'b100011111110;
		if(({row_reg, col_reg}>=18'b010111010010101000) && ({row_reg, col_reg}<18'b010111010010101010)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010111010010101010)) color_data = 12'b010010101011;
		if(({row_reg, col_reg}==18'b010111010010101011)) color_data = 12'b001010001010;
		if(({row_reg, col_reg}==18'b010111010010101100)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b010111010010101101)) color_data = 12'b001010011011;
		if(({row_reg, col_reg}==18'b010111010010101110)) color_data = 12'b001010011010;
		if(({row_reg, col_reg}==18'b010111010010101111)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010111010010110000)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010111010010110001) && ({row_reg, col_reg}<18'b010111010010110011)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010111010010110011) && ({row_reg, col_reg}<18'b010111010010110101)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010111010010110101) && ({row_reg, col_reg}<18'b010111010010110111)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010111010010110111)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010111010010111000)) color_data = 12'b011010111111;
		if(({row_reg, col_reg}==18'b010111010010111001)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010111010010111010)) color_data = 12'b001010001101;
		if(({row_reg, col_reg}==18'b010111010010111011)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111010010111100)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010111010010111101)) color_data = 12'b011011001111;
		if(({row_reg, col_reg}==18'b010111010010111110)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010111010010111111)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}>=18'b010111010011000000) && ({row_reg, col_reg}<18'b010111010011000010)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010111010011000010) && ({row_reg, col_reg}<18'b010111010011000111)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010111010011000111)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}>=18'b010111010011001000) && ({row_reg, col_reg}<18'b010111010011001010)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010111010011001010)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b010111010011001011)) color_data = 12'b011011001111;
		if(({row_reg, col_reg}==18'b010111010011001100)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010111010011001101)) color_data = 12'b001010001101;
		if(({row_reg, col_reg}==18'b010111010011001110)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}==18'b010111010011001111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111010011010000)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b010111010011010001) && ({row_reg, col_reg}<18'b010111010011010100)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010111010011010100) && ({row_reg, col_reg}<18'b010111010011011011)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}>=18'b010111010011011011) && ({row_reg, col_reg}<18'b010111010011011101)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111010011011101)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010111010011011110)) color_data = 12'b010110101110;
		if(({row_reg, col_reg}==18'b010111010011011111)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010111010011100000)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010111010011100001) && ({row_reg, col_reg}<18'b010111010011100011)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010111010011100011) && ({row_reg, col_reg}<18'b010111010011101000)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010111010011101000)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}>=18'b010111010011101001) && ({row_reg, col_reg}<18'b010111010011101110)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010111010011101110)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010111010011101111)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}>=18'b010111010011110000) && ({row_reg, col_reg}<18'b010111010011110101)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010111010011110101) && ({row_reg, col_reg}<18'b010111010011111000)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}>=18'b010111010011111000) && ({row_reg, col_reg}<18'b010111010011111101)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010111010011111101) && ({row_reg, col_reg}<18'b010111010100000000)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010111010100000000)) color_data = 12'b011110111111;
		if(({row_reg, col_reg}>=18'b010111010100000001) && ({row_reg, col_reg}<18'b010111010100000011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010111010100000011)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b010111010100000100)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}>=18'b010111010100000101) && ({row_reg, col_reg}<18'b010111010100001000)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010111010100001000)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b010111010100001001)) color_data = 12'b010010011101;
		if(({row_reg, col_reg}==18'b010111010100001010)) color_data = 12'b011010111111;
		if(({row_reg, col_reg}>=18'b010111010100001011) && ({row_reg, col_reg}<18'b010111010100001101)) color_data = 12'b011110111111;
		if(({row_reg, col_reg}==18'b010111010100001101)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b010111010100001110) && ({row_reg, col_reg}<18'b010111011000010000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010111011000010000) && ({row_reg, col_reg}<18'b010111011000010100)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b010111011000010100) && ({row_reg, col_reg}<18'b010111011000010110)) color_data = 12'b010110101111;
		if(({row_reg, col_reg}==18'b010111011000010110)) color_data = 12'b010010001110;
		if(({row_reg, col_reg}==18'b010111011000010111)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010111011000011000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010111011000011001) && ({row_reg, col_reg}<18'b010111011000011110)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010111011000011110)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010111011000011111)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b010111011000100000) && ({row_reg, col_reg}<18'b010111011000100011)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010111011000100011) && ({row_reg, col_reg}<18'b010111011000100101)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}>=18'b010111011000100101) && ({row_reg, col_reg}<18'b010111011000101001)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010111011000101001) && ({row_reg, col_reg}<18'b010111011000101011)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}>=18'b010111011000101011) && ({row_reg, col_reg}<18'b010111011000101101)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b010111011000101101) && ({row_reg, col_reg}<18'b010111011000101111)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010111011000101111)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}>=18'b010111011000110000) && ({row_reg, col_reg}<18'b010111011000110010)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}>=18'b010111011000110010) && ({row_reg, col_reg}<18'b010111011000110100)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b010111011000110100) && ({row_reg, col_reg}<18'b010111011000110110)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010111011000110110)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010111011000110111)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}==18'b010111011000111000)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}>=18'b010111011000111001) && ({row_reg, col_reg}<18'b010111011000111011)) color_data = 12'b011011001101;
		if(({row_reg, col_reg}==18'b010111011000111011)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}==18'b010111011000111100)) color_data = 12'b011011001110;
		if(({row_reg, col_reg}==18'b010111011000111101)) color_data = 12'b011111101111;
		if(({row_reg, col_reg}>=18'b010111011000111110) && ({row_reg, col_reg}<18'b010111011001000000)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}==18'b010111011001000000)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}>=18'b010111011001000001) && ({row_reg, col_reg}<18'b010111011001001000)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}>=18'b010111011001001000) && ({row_reg, col_reg}<18'b010111011001001010)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010111011001001010)) color_data = 12'b011111101111;
		if(({row_reg, col_reg}>=18'b010111011001001011) && ({row_reg, col_reg}<18'b010111011001010000)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}>=18'b010111011001010000) && ({row_reg, col_reg}<18'b010111011001010010)) color_data = 12'b011111011110;
		if(({row_reg, col_reg}==18'b010111011001010010)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}==18'b010111011001010011)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}>=18'b010111011001010100) && ({row_reg, col_reg}<18'b010111011001011000)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}==18'b010111011001011000)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010111011001011001)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010111011001011010) && ({row_reg, col_reg}<18'b010111011001011100)) color_data = 12'b100011111110;
		if(({row_reg, col_reg}==18'b010111011001011100)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010111011001011101)) color_data = 12'b100011101110;
		if(({row_reg, col_reg}==18'b010111011001011110)) color_data = 12'b010010011010;
		if(({row_reg, col_reg}==18'b010111011001011111)) color_data = 12'b010010001010;
		if(({row_reg, col_reg}==18'b010111011001100000)) color_data = 12'b011001111010;
		if(({row_reg, col_reg}==18'b010111011001100001)) color_data = 12'b011001101010;
		if(({row_reg, col_reg}==18'b010111011001100010)) color_data = 12'b011101111001;
		if(({row_reg, col_reg}>=18'b010111011001100011) && ({row_reg, col_reg}<18'b010111011001100101)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==18'b010111011001100101)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}>=18'b010111011001100110) && ({row_reg, col_reg}<18'b010111011001101000)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010111011001101000)) color_data = 12'b100001110110;
		if(({row_reg, col_reg}>=18'b010111011001101001) && ({row_reg, col_reg}<18'b010111011001101110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010111011001101110)) color_data = 12'b100001100110;
		if(({row_reg, col_reg}==18'b010111011001101111)) color_data = 12'b100001100101;
		if(({row_reg, col_reg}>=18'b010111011001110000) && ({row_reg, col_reg}<18'b010111011001110010)) color_data = 12'b100001100110;
		if(({row_reg, col_reg}>=18'b010111011001110010) && ({row_reg, col_reg}<18'b010111011001110100)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010111011001110100)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}==18'b010111011001110101)) color_data = 12'b011001101000;
		if(({row_reg, col_reg}==18'b010111011001110110)) color_data = 12'b011001101001;
		if(({row_reg, col_reg}==18'b010111011001110111)) color_data = 12'b011001111010;
		if(({row_reg, col_reg}==18'b010111011001111000)) color_data = 12'b010101111010;
		if(({row_reg, col_reg}==18'b010111011001111001)) color_data = 12'b001101111010;
		if(({row_reg, col_reg}==18'b010111011001111010)) color_data = 12'b010110101100;
		if(({row_reg, col_reg}==18'b010111011001111011)) color_data = 12'b100011011111;
		if(({row_reg, col_reg}>=18'b010111011001111100) && ({row_reg, col_reg}<18'b010111011001111111)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}==18'b010111011001111111)) color_data = 12'b010010101101;
		if(({row_reg, col_reg}==18'b010111011010000000)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b010111011010000001) && ({row_reg, col_reg}<18'b010111011010000100)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}>=18'b010111011010000100) && ({row_reg, col_reg}<18'b010111011010001000)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010111011010001000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010111011010001001) && ({row_reg, col_reg}<18'b010111011010001011)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b010111011010001011)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111011010001100)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b010111011010001101)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b010111011010001110)) color_data = 12'b010010011101;
		if(({row_reg, col_reg}>=18'b010111011010001111) && ({row_reg, col_reg}<18'b010111011010010010)) color_data = 12'b010010011100;
		if(({row_reg, col_reg}==18'b010111011010010010)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b010111011010010011)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010111011010010100)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010111011010010101) && ({row_reg, col_reg}<18'b010111011010011001)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010111011010011001)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111011010011010)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010111011010011011)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}>=18'b010111011010011100) && ({row_reg, col_reg}<18'b010111011010011110)) color_data = 12'b010010011101;
		if(({row_reg, col_reg}==18'b010111011010011110)) color_data = 12'b010010101101;
		if(({row_reg, col_reg}==18'b010111011010011111)) color_data = 12'b001110011011;
		if(({row_reg, col_reg}==18'b010111011010100000)) color_data = 12'b010110111100;
		if(({row_reg, col_reg}==18'b010111011010100001)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010111011010100010) && ({row_reg, col_reg}<18'b010111011010101011)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010111011010101011) && ({row_reg, col_reg}<18'b010111011010101101)) color_data = 12'b011111011110;
		if(({row_reg, col_reg}==18'b010111011010101101)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}>=18'b010111011010101110) && ({row_reg, col_reg}<18'b010111011010110000)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}>=18'b010111011010110000) && ({row_reg, col_reg}<18'b010111011010110011)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010111011010110011)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010111011010110100)) color_data = 12'b001110011010;
		if(({row_reg, col_reg}==18'b010111011010110101)) color_data = 12'b001110011011;
		if(({row_reg, col_reg}==18'b010111011010110110)) color_data = 12'b010010101101;
		if(({row_reg, col_reg}==18'b010111011010110111)) color_data = 12'b001110011100;
		if(({row_reg, col_reg}==18'b010111011010111000)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}>=18'b010111011010111001) && ({row_reg, col_reg}<18'b010111011010111100)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111011010111100)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b010111011010111101) && ({row_reg, col_reg}<18'b010111011010111111)) color_data = 12'b010010011101;
		if(({row_reg, col_reg}==18'b010111011010111111)) color_data = 12'b010010011100;
		if(({row_reg, col_reg}>=18'b010111011011000000) && ({row_reg, col_reg}<18'b010111011011000010)) color_data = 12'b010010101100;
		if(({row_reg, col_reg}==18'b010111011011000010)) color_data = 12'b001110101100;
		if(({row_reg, col_reg}>=18'b010111011011000011) && ({row_reg, col_reg}<18'b010111011011000101)) color_data = 12'b001110011100;
		if(({row_reg, col_reg}>=18'b010111011011000101) && ({row_reg, col_reg}<18'b010111011011000111)) color_data = 12'b001110101100;
		if(({row_reg, col_reg}>=18'b010111011011000111) && ({row_reg, col_reg}<18'b010111011011001001)) color_data = 12'b001110011100;
		if(({row_reg, col_reg}==18'b010111011011001001)) color_data = 12'b010010101101;
		if(({row_reg, col_reg}==18'b010111011011001010)) color_data = 12'b001110011101;
		if(({row_reg, col_reg}==18'b010111011011001011)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b010111011011001100)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010111011011001101)) color_data = 12'b001010001101;
		if(({row_reg, col_reg}>=18'b010111011011001110) && ({row_reg, col_reg}<18'b010111011011010011)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010111011011010011) && ({row_reg, col_reg}<18'b010111011011011011)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b010111011011011011)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010111011011011100)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010111011011011101)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111011011011110)) color_data = 12'b010010011110;
		if(({row_reg, col_reg}==18'b010111011011011111)) color_data = 12'b011010111111;
		if(({row_reg, col_reg}==18'b010111011011100000)) color_data = 12'b011110111110;
		if(({row_reg, col_reg}==18'b010111011011100001)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}>=18'b010111011011100010) && ({row_reg, col_reg}<18'b010111011011100110)) color_data = 12'b011110111110;
		if(({row_reg, col_reg}>=18'b010111011011100110) && ({row_reg, col_reg}<18'b010111011011101000)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==18'b010111011011101000)) color_data = 12'b011110111110;
		if(({row_reg, col_reg}>=18'b010111011011101001) && ({row_reg, col_reg}<18'b010111011011101011)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==18'b010111011011101011)) color_data = 12'b011011001110;
		if(({row_reg, col_reg}==18'b010111011011101100)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==18'b010111011011101101)) color_data = 12'b010010101101;
		if(({row_reg, col_reg}==18'b010111011011101110)) color_data = 12'b001110011100;
		if(({row_reg, col_reg}==18'b010111011011101111)) color_data = 12'b010010101101;
		if(({row_reg, col_reg}==18'b010111011011110000)) color_data = 12'b001110011100;
		if(({row_reg, col_reg}==18'b010111011011110001)) color_data = 12'b010010101100;
		if(({row_reg, col_reg}>=18'b010111011011110010) && ({row_reg, col_reg}<18'b010111011011110100)) color_data = 12'b001110011100;
		if(({row_reg, col_reg}==18'b010111011011110100)) color_data = 12'b010010011100;
		if(({row_reg, col_reg}==18'b010111011011110101)) color_data = 12'b010010011101;
		if(({row_reg, col_reg}==18'b010111011011110110)) color_data = 12'b010010011110;
		if(({row_reg, col_reg}>=18'b010111011011110111) && ({row_reg, col_reg}<18'b010111011011111001)) color_data = 12'b010010011101;
		if(({row_reg, col_reg}==18'b010111011011111001)) color_data = 12'b001110011100;
		if(({row_reg, col_reg}==18'b010111011011111010)) color_data = 12'b010010101100;
		if(({row_reg, col_reg}==18'b010111011011111011)) color_data = 12'b001110101100;
		if(({row_reg, col_reg}>=18'b010111011011111100) && ({row_reg, col_reg}<18'b010111011011111110)) color_data = 12'b010010101101;
		if(({row_reg, col_reg}>=18'b010111011011111110) && ({row_reg, col_reg}<18'b010111011100000000)) color_data = 12'b010010011100;
		if(({row_reg, col_reg}>=18'b010111011100000000) && ({row_reg, col_reg}<18'b010111011100000101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010111011100000101) && ({row_reg, col_reg}<18'b010111011100000111)) color_data = 12'b011010011110;
		if(({row_reg, col_reg}==18'b010111011100000111)) color_data = 12'b010110101110;
		if(({row_reg, col_reg}>=18'b010111011100001000) && ({row_reg, col_reg}<18'b010111011100001010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010111011100001010)) color_data = 12'b011010101111;

		if(({row_reg, col_reg}>=18'b010111011100001011) && ({row_reg, col_reg}<18'b010111100000010000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010111100000010000) && ({row_reg, col_reg}<18'b010111100000010110)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b010111100000010110)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}>=18'b010111100000010111) && ({row_reg, col_reg}<18'b010111100000100000)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b010111100000100000) && ({row_reg, col_reg}<18'b010111100000100101)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111100000100101)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010111100000100110)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010111100000100111)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b010111100000101000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010111100000101001) && ({row_reg, col_reg}<18'b010111100000101100)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}>=18'b010111100000101100) && ({row_reg, col_reg}<18'b010111100000101110)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010111100000101110) && ({row_reg, col_reg}<18'b010111100000110000)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b010111100000110000) && ({row_reg, col_reg}<18'b010111100000110011)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010111100000110011)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010111100000110100)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b010111100000110101) && ({row_reg, col_reg}<18'b010111100000110111)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010111100000110111)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b010111100000111000)) color_data = 12'b010110101101;
		if(({row_reg, col_reg}==18'b010111100000111001)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}>=18'b010111100000111010) && ({row_reg, col_reg}<18'b010111100000111100)) color_data = 12'b010110111100;
		if(({row_reg, col_reg}==18'b010111100000111100)) color_data = 12'b011111001110;
		if(({row_reg, col_reg}==18'b010111100000111101)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010111100000111110) && ({row_reg, col_reg}<18'b010111100001000000)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010111100001000000) && ({row_reg, col_reg}<18'b010111100001001001)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010111100001001001) && ({row_reg, col_reg}<18'b010111100001010000)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010111100001010000) && ({row_reg, col_reg}<18'b010111100001010110)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010111100001010110) && ({row_reg, col_reg}<18'b010111100001011000)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010111100001011000)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010111100001011001)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010111100001011010)) color_data = 12'b100011111110;
		if(({row_reg, col_reg}==18'b010111100001011011)) color_data = 12'b011111111110;
		if(({row_reg, col_reg}==18'b010111100001011100)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010111100001011101)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010111100001011110)) color_data = 12'b001110001011;
		if(({row_reg, col_reg}==18'b010111100001011111)) color_data = 12'b001101111010;
		if(({row_reg, col_reg}==18'b010111100001100000)) color_data = 12'b010101111011;
		if(({row_reg, col_reg}==18'b010111100001100001)) color_data = 12'b010101101010;
		if(({row_reg, col_reg}==18'b010111100001100010)) color_data = 12'b011001101001;
		if(({row_reg, col_reg}==18'b010111100001100011)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}==18'b010111100001100100)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010111100001100101)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}==18'b010111100001100110)) color_data = 12'b011001100101;
		if(({row_reg, col_reg}==18'b010111100001100111)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010111100001101000) && ({row_reg, col_reg}<18'b010111100001101010)) color_data = 12'b011101100111;
		if(({row_reg, col_reg}>=18'b010111100001101010) && ({row_reg, col_reg}<18'b010111100001101100)) color_data = 12'b011101110111;
		if(({row_reg, col_reg}>=18'b010111100001101100) && ({row_reg, col_reg}<18'b010111100001101110)) color_data = 12'b011101100110;
		if(({row_reg, col_reg}>=18'b010111100001101110) && ({row_reg, col_reg}<18'b010111100001110001)) color_data = 12'b011101100101;
		if(({row_reg, col_reg}>=18'b010111100001110001) && ({row_reg, col_reg}<18'b010111100001110011)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010111100001110011)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}==18'b010111100001110100)) color_data = 12'b011001111000;
		if(({row_reg, col_reg}>=18'b010111100001110101) && ({row_reg, col_reg}<18'b010111100001110111)) color_data = 12'b010101101001;
		if(({row_reg, col_reg}==18'b010111100001110111)) color_data = 12'b010101111011;
		if(({row_reg, col_reg}==18'b010111100001111000)) color_data = 12'b010001111011;
		if(({row_reg, col_reg}==18'b010111100001111001)) color_data = 12'b001101111010;
		if(({row_reg, col_reg}==18'b010111100001111010)) color_data = 12'b010110101101;
		if(({row_reg, col_reg}>=18'b010111100001111011) && ({row_reg, col_reg}<18'b010111100001111111)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010111100001111111)) color_data = 12'b010110111101;
		if(({row_reg, col_reg}>=18'b010111100010000000) && ({row_reg, col_reg}<18'b010111100010000010)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b010111100010000010) && ({row_reg, col_reg}<18'b010111100010000100)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}>=18'b010111100010000100) && ({row_reg, col_reg}<18'b010111100010001000)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010111100010001000)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010111100010001001)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111100010001010)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}>=18'b010111100010001011) && ({row_reg, col_reg}<18'b010111100010001101)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010111100010001101) && ({row_reg, col_reg}<18'b010111100010001111)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b010111100010001111)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b010111100010010000)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}>=18'b010111100010010001) && ({row_reg, col_reg}<18'b010111100010010011)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b010111100010010011) && ({row_reg, col_reg}<18'b010111100010011001)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111100010011001)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b010111100010011010) && ({row_reg, col_reg}<18'b010111100010011100)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111100010011100)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010111100010011101)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b010111100010011110)) color_data = 12'b001110001011;
		if(({row_reg, col_reg}==18'b010111100010011111)) color_data = 12'b001001111010;
		if(({row_reg, col_reg}==18'b010111100010100000)) color_data = 12'b010010101011;
		if(({row_reg, col_reg}==18'b010111100010100001)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010111100010100010) && ({row_reg, col_reg}<18'b010111100010100110)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010111100010100110)) color_data = 12'b100011111110;
		if(({row_reg, col_reg}>=18'b010111100010100111) && ({row_reg, col_reg}<18'b010111100010101011)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010111100010101011) && ({row_reg, col_reg}<18'b010111100010101110)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010111100010101110)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010111100010101111) && ({row_reg, col_reg}<18'b010111100010110011)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010111100010110011)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}==18'b010111100010110100)) color_data = 12'b001001111010;
		if(({row_reg, col_reg}==18'b010111100010110101)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b010111100010110110)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b010111100010110111)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010111100010111000)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}==18'b010111100010111001)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111100010111010)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b010111100010111011)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010111100010111100)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010111100010111101) && ({row_reg, col_reg}<18'b010111100011000000)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b010111100011000000) && ({row_reg, col_reg}<18'b010111100011000011)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b010111100011000011)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b010111100011000100)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b010111100011000101)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b010111100011000110)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b010111100011000111)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}>=18'b010111100011001000) && ({row_reg, col_reg}<18'b010111100011001011)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010111100011001011)) color_data = 12'b001010001101;
		if(({row_reg, col_reg}>=18'b010111100011001100) && ({row_reg, col_reg}<18'b010111100011010000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010111100011010000) && ({row_reg, col_reg}<18'b010111100011011011)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b010111100011011011)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010111100011011100)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010111100011011101)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010111100011011110)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}==18'b010111100011011111)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b010111100011100000) && ({row_reg, col_reg}<18'b010111100011100111)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}>=18'b010111100011100111) && ({row_reg, col_reg}<18'b010111100011101001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010111100011101001)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==18'b010111100011101010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010111100011101011) && ({row_reg, col_reg}<18'b010111100011101101)) color_data = 12'b010110101110;
		if(({row_reg, col_reg}==18'b010111100011101101)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b010111100011101110)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010111100011101111)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b010111100011110000)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b010111100011110001) && ({row_reg, col_reg}<18'b010111100011110100)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b010111100011110100)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b010111100011110101) && ({row_reg, col_reg}<18'b010111100011110111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111100011110111)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010111100011111000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111100011111001)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010111100011111010)) color_data = 12'b000101111100;
		if(({row_reg, col_reg}==18'b010111100011111011)) color_data = 12'b000101111011;
		if(({row_reg, col_reg}>=18'b010111100011111100) && ({row_reg, col_reg}<18'b010111100011111110)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010111100011111110)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b010111100011111111)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b010111100100000000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010111100100000001)) color_data = 12'b011110111111;
		if(({row_reg, col_reg}>=18'b010111100100000010) && ({row_reg, col_reg}<18'b010111100100000110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010111100100000110) && ({row_reg, col_reg}<18'b010111100100001010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010111100100001010)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b010111100100001011) && ({row_reg, col_reg}<18'b010111100100001101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010111100100001101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b010111100100001110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010111100100001111)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b010111100100010000) && ({row_reg, col_reg}<18'b010111101000010011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010111101000010011) && ({row_reg, col_reg}<18'b010111101000010110)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b010111101000010110)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==18'b010111101000010111)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010111101000011000)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}>=18'b010111101000011001) && ({row_reg, col_reg}<18'b010111101000100011)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b010111101000100011) && ({row_reg, col_reg}<18'b010111101000100110)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111101000100110)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010111101000100111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010111101000101000) && ({row_reg, col_reg}<18'b010111101000101100)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}>=18'b010111101000101100) && ({row_reg, col_reg}<18'b010111101000101110)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b010111101000101110) && ({row_reg, col_reg}<18'b010111101000110001)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010111101000110001)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}>=18'b010111101000110010) && ({row_reg, col_reg}<18'b010111101000110111)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010111101000110111)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}==18'b010111101000111000)) color_data = 12'b010110101110;
		if(({row_reg, col_reg}==18'b010111101000111001)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==18'b010111101000111010)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}==18'b010111101000111011)) color_data = 12'b010110111100;
		if(({row_reg, col_reg}==18'b010111101000111100)) color_data = 12'b011111011110;
		if(({row_reg, col_reg}>=18'b010111101000111101) && ({row_reg, col_reg}<18'b010111101001000000)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010111101001000000) && ({row_reg, col_reg}<18'b010111101001001000)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010111101001001000)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010111101001001001) && ({row_reg, col_reg}<18'b010111101001010111)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010111101001010111)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010111101001011000) && ({row_reg, col_reg}<18'b010111101001011010)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010111101001011010)) color_data = 12'b100011111110;
		if(({row_reg, col_reg}==18'b010111101001011011)) color_data = 12'b011111111110;
		if(({row_reg, col_reg}==18'b010111101001011100)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010111101001011101)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010111101001011110)) color_data = 12'b010010011100;
		if(({row_reg, col_reg}==18'b010111101001011111)) color_data = 12'b001001111010;
		if(({row_reg, col_reg}==18'b010111101001100000)) color_data = 12'b010001111011;
		if(({row_reg, col_reg}==18'b010111101001100001)) color_data = 12'b010101111011;
		if(({row_reg, col_reg}==18'b010111101001100010)) color_data = 12'b010101111010;
		if(({row_reg, col_reg}==18'b010111101001100011)) color_data = 12'b011001111001;
		if(({row_reg, col_reg}==18'b010111101001100100)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==18'b010111101001100101)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}==18'b010111101001100110)) color_data = 12'b011001100110;
		if(({row_reg, col_reg}==18'b010111101001100111)) color_data = 12'b011001110111;
		if(({row_reg, col_reg}==18'b010111101001101000)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}==18'b010111101001101001)) color_data = 12'b011001101000;
		if(({row_reg, col_reg}>=18'b010111101001101010) && ({row_reg, col_reg}<18'b010111101001101101)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}>=18'b010111101001101101) && ({row_reg, col_reg}<18'b010111101001110001)) color_data = 12'b011101110110;
		if(({row_reg, col_reg}==18'b010111101001110001)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}==18'b010111101001110010)) color_data = 12'b011001100111;
		if(({row_reg, col_reg}==18'b010111101001110011)) color_data = 12'b010101101000;
		if(({row_reg, col_reg}==18'b010111101001110100)) color_data = 12'b010101111001;
		if(({row_reg, col_reg}==18'b010111101001110101)) color_data = 12'b010101111010;
		if(({row_reg, col_reg}==18'b010111101001110110)) color_data = 12'b010001101010;
		if(({row_reg, col_reg}==18'b010111101001110111)) color_data = 12'b010001111011;
		if(({row_reg, col_reg}>=18'b010111101001111000) && ({row_reg, col_reg}<18'b010111101001111010)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010111101001111010)) color_data = 12'b010110101101;
		if(({row_reg, col_reg}==18'b010111101001111011)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}>=18'b010111101001111100) && ({row_reg, col_reg}<18'b010111101001111110)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010111101001111110)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010111101001111111)) color_data = 12'b010110111101;
		if(({row_reg, col_reg}==18'b010111101010000000)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010111101010000001)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b010111101010000010)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}>=18'b010111101010000011) && ({row_reg, col_reg}<18'b010111101010000111)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b010111101010000111) && ({row_reg, col_reg}<18'b010111101010001001)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010111101010001001)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010111101010001010) && ({row_reg, col_reg}<18'b010111101010001101)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b010111101010001101) && ({row_reg, col_reg}<18'b010111101010010001)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111101010010001)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b010111101010010010) && ({row_reg, col_reg}<18'b010111101010010111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010111101010010111) && ({row_reg, col_reg}<18'b010111101010011001)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010111101010011001)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}>=18'b010111101010011010) && ({row_reg, col_reg}<18'b010111101010011100)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010111101010011100)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}==18'b010111101010011101)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010111101010011110)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b010111101010011111)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b010111101010100000)) color_data = 12'b010010101100;
		if(({row_reg, col_reg}==18'b010111101010100001)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010111101010100010)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010111101010100011) && ({row_reg, col_reg}<18'b010111101010101101)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010111101010101101)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010111101010101110) && ({row_reg, col_reg}<18'b010111101010110001)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010111101010110001) && ({row_reg, col_reg}<18'b010111101010110011)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010111101010110011)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}==18'b010111101010110100)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b010111101010110101)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b010111101010110110)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010111101010110111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111101010111000)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}==18'b010111101010111001)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}>=18'b010111101010111010) && ({row_reg, col_reg}<18'b010111101010111110)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b010111101010111110) && ({row_reg, col_reg}<18'b010111101011000000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010111101011000000) && ({row_reg, col_reg}<18'b010111101011000101)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010111101011000101)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010111101011000110)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b010111101011000111)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010111101011001000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111101011001001)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}>=18'b010111101011001010) && ({row_reg, col_reg}<18'b010111101011001100)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111101011001100)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}>=18'b010111101011001101) && ({row_reg, col_reg}<18'b010111101011010000)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b010111101011010000) && ({row_reg, col_reg}<18'b010111101011011100)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b010111101011011100) && ({row_reg, col_reg}<18'b010111101011011110)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010111101011011110)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}==18'b010111101011011111)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b010111101011100000)) color_data = 12'b011110111110;
		if(({row_reg, col_reg}==18'b010111101011100001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010111101011100010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010111101011100011) && ({row_reg, col_reg}<18'b010111101011100110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010111101011100110)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}>=18'b010111101011100111) && ({row_reg, col_reg}<18'b010111101011101011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010111101011101011)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b010111101011101100)) color_data = 12'b010110101111;
		if(({row_reg, col_reg}==18'b010111101011101101)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b010111101011101110)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111101011101111)) color_data = 12'b001010001110;
		if(({row_reg, col_reg}==18'b010111101011110000)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010111101011110001)) color_data = 12'b001010001101;
		if(({row_reg, col_reg}==18'b010111101011110010)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010111101011110011)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}>=18'b010111101011110100) && ({row_reg, col_reg}<18'b010111101011110110)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b010111101011110110) && ({row_reg, col_reg}<18'b010111101011111001)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010111101011111001)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b010111101011111010) && ({row_reg, col_reg}<18'b010111101011111100)) color_data = 12'b001010001101;
		if(({row_reg, col_reg}==18'b010111101011111100)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}==18'b010111101011111101)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010111101011111110)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010111101011111111)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}==18'b010111101100000000)) color_data = 12'b010110011101;
		if(({row_reg, col_reg}==18'b010111101100000001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010111101100000010) && ({row_reg, col_reg}<18'b010111101100000101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b010111101100000101)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b010111101100000110)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}>=18'b010111101100000111) && ({row_reg, col_reg}<18'b010111101100001010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010111101100001010)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}>=18'b010111101100001011) && ({row_reg, col_reg}<18'b010111101100001111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010111101100001111)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b010111101100010000) && ({row_reg, col_reg}<18'b010111110000010101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010111110000010101)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b010111110000010110)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}>=18'b010111110000010111) && ({row_reg, col_reg}<18'b010111110000011010)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}>=18'b010111110000011010) && ({row_reg, col_reg}<18'b010111110000011101)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010111110000011101)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111110000011110)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b010111110000011111) && ({row_reg, col_reg}<18'b010111110000100010)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010111110000100010) && ({row_reg, col_reg}<18'b010111110000100101)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b010111110000100101) && ({row_reg, col_reg}<18'b010111110000101000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010111110000101000) && ({row_reg, col_reg}<18'b010111110000101100)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}>=18'b010111110000101100) && ({row_reg, col_reg}<18'b010111110000101110)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010111110000101110) && ({row_reg, col_reg}<18'b010111110000110000)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010111110000110000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111110000110001)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010111110000110010)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b010111110000110011) && ({row_reg, col_reg}<18'b010111110000110111)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010111110000110111)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b010111110000111000)) color_data = 12'b010110101110;
		if(({row_reg, col_reg}==18'b010111110000111001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010111110000111010)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==18'b010111110000111011)) color_data = 12'b010110101100;
		if(({row_reg, col_reg}==18'b010111110000111100)) color_data = 12'b011111001110;
		if(({row_reg, col_reg}==18'b010111110000111101)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}>=18'b010111110000111110) && ({row_reg, col_reg}<18'b010111110001000001)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010111110001000001)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010111110001000010) && ({row_reg, col_reg}<18'b010111110001000100)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010111110001000100) && ({row_reg, col_reg}<18'b010111110001000110)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010111110001000110) && ({row_reg, col_reg}<18'b010111110001001000)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010111110001001000) && ({row_reg, col_reg}<18'b010111110001010001)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010111110001010001)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010111110001010010) && ({row_reg, col_reg}<18'b010111110001010101)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010111110001010101) && ({row_reg, col_reg}<18'b010111110001011010)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b010111110001011010) && ({row_reg, col_reg}<18'b010111110001011101)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010111110001011101)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010111110001011110)) color_data = 12'b001110011100;
		if(({row_reg, col_reg}==18'b010111110001011111)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b010111110001100000)) color_data = 12'b001001111010;
		if(({row_reg, col_reg}==18'b010111110001100001)) color_data = 12'b001101111010;
		if(({row_reg, col_reg}==18'b010111110001100010)) color_data = 12'b001101111001;
		if(({row_reg, col_reg}==18'b010111110001100011)) color_data = 12'b010001100111;
		if(({row_reg, col_reg}>=18'b010111110001100100) && ({row_reg, col_reg}<18'b010111110001100110)) color_data = 12'b010001100110;
		if(({row_reg, col_reg}>=18'b010111110001100110) && ({row_reg, col_reg}<18'b010111110001101000)) color_data = 12'b010101110111;
		if(({row_reg, col_reg}==18'b010111110001101000)) color_data = 12'b010101101000;
		if(({row_reg, col_reg}==18'b010111110001101001)) color_data = 12'b011001101001;
		if(({row_reg, col_reg}==18'b010111110001101010)) color_data = 12'b011001111001;
		if(({row_reg, col_reg}==18'b010111110001101011)) color_data = 12'b011001101000;
		if(({row_reg, col_reg}==18'b010111110001101100)) color_data = 12'b010101100111;
		if(({row_reg, col_reg}==18'b010111110001101101)) color_data = 12'b010101100110;
		if(({row_reg, col_reg}>=18'b010111110001101110) && ({row_reg, col_reg}<18'b010111110001110000)) color_data = 12'b010101100101;
		if(({row_reg, col_reg}==18'b010111110001110000)) color_data = 12'b011001110110;
		if(({row_reg, col_reg}==18'b010111110001110001)) color_data = 12'b010101100111;
		if(({row_reg, col_reg}==18'b010111110001110010)) color_data = 12'b010101111000;
		if(({row_reg, col_reg}==18'b010111110001110011)) color_data = 12'b010101111001;
		if(({row_reg, col_reg}>=18'b010111110001110100) && ({row_reg, col_reg}<18'b010111110001110110)) color_data = 12'b010001111010;
		if(({row_reg, col_reg}==18'b010111110001110110)) color_data = 12'b001101111011;
		if(({row_reg, col_reg}>=18'b010111110001110111) && ({row_reg, col_reg}<18'b010111110001111001)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010111110001111001)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b010111110001111010)) color_data = 12'b010110101110;
		if(({row_reg, col_reg}==18'b010111110001111011)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}>=18'b010111110001111100) && ({row_reg, col_reg}<18'b010111110001111110)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010111110001111110)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010111110001111111)) color_data = 12'b010110111110;
		if(({row_reg, col_reg}>=18'b010111110010000000) && ({row_reg, col_reg}<18'b010111110010000010)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b010111110010000010) && ({row_reg, col_reg}<18'b010111110010000100)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010111110010000100) && ({row_reg, col_reg}<18'b010111110010001001)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b010111110010001001) && ({row_reg, col_reg}<18'b010111110010001011)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b010111110010001011) && ({row_reg, col_reg}<18'b010111110010001101)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b010111110010001101) && ({row_reg, col_reg}<18'b010111110010010000)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}>=18'b010111110010010000) && ({row_reg, col_reg}<18'b010111110010010010)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010111110010010010)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}>=18'b010111110010010011) && ({row_reg, col_reg}<18'b010111110010010111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111110010010111)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010111110010011000)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}>=18'b010111110010011001) && ({row_reg, col_reg}<18'b010111110010011101)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b010111110010011101) && ({row_reg, col_reg}<18'b010111110010011111)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010111110010011111)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010111110010100000)) color_data = 12'b010110101101;
		if(({row_reg, col_reg}==18'b010111110010100001)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}>=18'b010111110010100010) && ({row_reg, col_reg}<18'b010111110010101010)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010111110010101010)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b010111110010101011) && ({row_reg, col_reg}<18'b010111110010110011)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b010111110010110011)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}==18'b010111110010110100)) color_data = 12'b001110011100;
		if(({row_reg, col_reg}==18'b010111110010110101)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b010111110010110110) && ({row_reg, col_reg}<18'b010111110010111000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111110010111000)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}>=18'b010111110010111001) && ({row_reg, col_reg}<18'b010111110011000000)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010111110011000000)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010111110011000001)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b010111110011000010) && ({row_reg, col_reg}<18'b010111110011000100)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010111110011000100)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}>=18'b010111110011000101) && ({row_reg, col_reg}<18'b010111110011000111)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b010111110011000111) && ({row_reg, col_reg}<18'b010111110011001001)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111110011001001)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}>=18'b010111110011001010) && ({row_reg, col_reg}<18'b010111110011001100)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010111110011001100) && ({row_reg, col_reg}<18'b010111110011001110)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010111110011001110)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b010111110011001111) && ({row_reg, col_reg}<18'b010111110011010001)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010111110011010001) && ({row_reg, col_reg}<18'b010111110011010011)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010111110011010011)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111110011010100)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b010111110011010101) && ({row_reg, col_reg}<18'b010111110011011001)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}>=18'b010111110011011001) && ({row_reg, col_reg}<18'b010111110011011101)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010111110011011101)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010111110011011110)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}>=18'b010111110011011111) && ({row_reg, col_reg}<18'b010111110011100111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010111110011100111)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010111110011101000) && ({row_reg, col_reg}<18'b010111110011101011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010111110011101011)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b010111110011101100)) color_data = 12'b010110101111;
		if(({row_reg, col_reg}==18'b010111110011101101)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b010111110011101110)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b010111110011101111) && ({row_reg, col_reg}<18'b010111110011110001)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111110011110001)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}>=18'b010111110011110010) && ({row_reg, col_reg}<18'b010111110011110101)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}>=18'b010111110011110101) && ({row_reg, col_reg}<18'b010111110011111000)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010111110011111000)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010111110011111001)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b010111110011111010) && ({row_reg, col_reg}<18'b010111110011111100)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111110011111100)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b010111110011111101)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010111110011111110)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010111110011111111)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}==18'b010111110100000000)) color_data = 12'b010110011101;
		if(({row_reg, col_reg}==18'b010111110100000001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010111110100000010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010111110100000011) && ({row_reg, col_reg}<18'b010111110100000110)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b010111110100000110)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}>=18'b010111110100000111) && ({row_reg, col_reg}<18'b010111110100001101)) color_data = 12'b011010101110;

		if(({row_reg, col_reg}>=18'b010111110100001101) && ({row_reg, col_reg}<18'b010111111000000000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010111111000000000) && ({row_reg, col_reg}<18'b010111111000010101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010111111000010101)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b010111111000010110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010111111000010111) && ({row_reg, col_reg}<18'b010111111000011001)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}>=18'b010111111000011001) && ({row_reg, col_reg}<18'b010111111000100101)) color_data = 12'b010010001110;
		if(({row_reg, col_reg}==18'b010111111000100101)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b010111111000100110) && ({row_reg, col_reg}<18'b010111111000101001)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010111111000101001) && ({row_reg, col_reg}<18'b010111111000101100)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b010111111000101100)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111111000101101)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010111111000101110)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}>=18'b010111111000101111) && ({row_reg, col_reg}<18'b010111111000110011)) color_data = 12'b010010001110;
		if(({row_reg, col_reg}>=18'b010111111000110011) && ({row_reg, col_reg}<18'b010111111000110111)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}==18'b010111111000110111)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==18'b010111111000111000)) color_data = 12'b010110101110;
		if(({row_reg, col_reg}==18'b010111111000111001)) color_data = 12'b011010111111;
		if(({row_reg, col_reg}==18'b010111111000111010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010111111000111011)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}==18'b010111111000111100)) color_data = 12'b011111001110;
		if(({row_reg, col_reg}>=18'b010111111000111101) && ({row_reg, col_reg}<18'b010111111001000000)) color_data = 12'b100011011111;
		if(({row_reg, col_reg}==18'b010111111001000000)) color_data = 12'b011111101111;
		if(({row_reg, col_reg}>=18'b010111111001000001) && ({row_reg, col_reg}<18'b010111111001000011)) color_data = 12'b011011011110;
		if(({row_reg, col_reg}==18'b010111111001000011)) color_data = 12'b011011011111;
		if(({row_reg, col_reg}>=18'b010111111001000100) && ({row_reg, col_reg}<18'b010111111001000110)) color_data = 12'b011011011110;
		if(({row_reg, col_reg}==18'b010111111001000110)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}>=18'b010111111001000111) && ({row_reg, col_reg}<18'b010111111001001111)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b010111111001001111)) color_data = 12'b011111111110;
		if(({row_reg, col_reg}==18'b010111111001010000)) color_data = 12'b011011001110;
		if(({row_reg, col_reg}==18'b010111111001010001)) color_data = 12'b011011011111;
		if(({row_reg, col_reg}>=18'b010111111001010010) && ({row_reg, col_reg}<18'b010111111001010100)) color_data = 12'b011011011110;
		if(({row_reg, col_reg}==18'b010111111001010100)) color_data = 12'b011011001110;
		if(({row_reg, col_reg}==18'b010111111001010101)) color_data = 12'b011011011110;
		if(({row_reg, col_reg}==18'b010111111001010110)) color_data = 12'b011011001110;
		if(({row_reg, col_reg}>=18'b010111111001010111) && ({row_reg, col_reg}<18'b010111111001011010)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}>=18'b010111111001011010) && ({row_reg, col_reg}<18'b010111111001011100)) color_data = 12'b011011011110;
		if(({row_reg, col_reg}>=18'b010111111001011100) && ({row_reg, col_reg}<18'b010111111001011110)) color_data = 12'b010111001110;
		if(({row_reg, col_reg}==18'b010111111001011110)) color_data = 12'b010110111110;
		if(({row_reg, col_reg}==18'b010111111001011111)) color_data = 12'b010110101110;
		if(({row_reg, col_reg}==18'b010111111001100000)) color_data = 12'b010010101101;
		if(({row_reg, col_reg}==18'b010111111001100001)) color_data = 12'b010110101100;
		if(({row_reg, col_reg}==18'b010111111001100010)) color_data = 12'b011010101011;
		if(({row_reg, col_reg}==18'b010111111001100011)) color_data = 12'b010110011010;
		if(({row_reg, col_reg}>=18'b010111111001100100) && ({row_reg, col_reg}<18'b010111111001100110)) color_data = 12'b011010011001;
		if(({row_reg, col_reg}==18'b010111111001100110)) color_data = 12'b011110101001;
		if(({row_reg, col_reg}==18'b010111111001100111)) color_data = 12'b011010011001;
		if(({row_reg, col_reg}==18'b010111111001101000)) color_data = 12'b010101101000;
		if(({row_reg, col_reg}==18'b010111111001101001)) color_data = 12'b010101111001;
		if(({row_reg, col_reg}==18'b010111111001101010)) color_data = 12'b011001111001;
		if(({row_reg, col_reg}==18'b010111111001101011)) color_data = 12'b010101111001;
		if(({row_reg, col_reg}==18'b010111111001101100)) color_data = 12'b011010001001;
		if(({row_reg, col_reg}==18'b010111111001101101)) color_data = 12'b011110011001;
		if(({row_reg, col_reg}>=18'b010111111001101110) && ({row_reg, col_reg}<18'b010111111001110000)) color_data = 12'b011110011000;
		if(({row_reg, col_reg}==18'b010111111001110000)) color_data = 12'b011110001001;
		if(({row_reg, col_reg}==18'b010111111001110001)) color_data = 12'b010101111000;
		if(({row_reg, col_reg}==18'b010111111001110010)) color_data = 12'b010101111001;
		if(({row_reg, col_reg}>=18'b010111111001110011) && ({row_reg, col_reg}<18'b010111111001110101)) color_data = 12'b010001111010;
		if(({row_reg, col_reg}==18'b010111111001110101)) color_data = 12'b010010001100;
		if(({row_reg, col_reg}>=18'b010111111001110110) && ({row_reg, col_reg}<18'b010111111001111000)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010111111001111000)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010111111001111001)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b010111111001111010)) color_data = 12'b010010011101;
		if(({row_reg, col_reg}==18'b010111111001111011)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}==18'b010111111001111100)) color_data = 12'b011011011110;
		if(({row_reg, col_reg}>=18'b010111111001111101) && ({row_reg, col_reg}<18'b010111111001111111)) color_data = 12'b011011001110;
		if(({row_reg, col_reg}==18'b010111111001111111)) color_data = 12'b010010101101;
		if(({row_reg, col_reg}==18'b010111111010000000)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}>=18'b010111111010000001) && ({row_reg, col_reg}<18'b010111111010000011)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010111111010000011) && ({row_reg, col_reg}<18'b010111111010000111)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}>=18'b010111111010000111) && ({row_reg, col_reg}<18'b010111111010001010)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010111111010001010)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010111111010001011)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111111010001100)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010111111010001101)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b010111111010001110) && ({row_reg, col_reg}<18'b010111111010010000)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b010111111010010000)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010111111010010001)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b010111111010010010) && ({row_reg, col_reg}<18'b010111111010010100)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b010111111010010100) && ({row_reg, col_reg}<18'b010111111010010111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010111111010010111) && ({row_reg, col_reg}<18'b010111111010011101)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b010111111010011101) && ({row_reg, col_reg}<18'b010111111010011111)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010111111010011111)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b010111111010100000)) color_data = 12'b010010011100;
		if(({row_reg, col_reg}==18'b010111111010100001)) color_data = 12'b011011001111;
		if(({row_reg, col_reg}>=18'b010111111010100010) && ({row_reg, col_reg}<18'b010111111010100100)) color_data = 12'b011011001110;
		if(({row_reg, col_reg}==18'b010111111010100100)) color_data = 12'b011011001101;
		if(({row_reg, col_reg}==18'b010111111010100101)) color_data = 12'b011111011110;
		if(({row_reg, col_reg}==18'b010111111010100110)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b010111111010100111)) color_data = 12'b011111011110;
		if(({row_reg, col_reg}==18'b010111111010101000)) color_data = 12'b011111101111;
		if(({row_reg, col_reg}>=18'b010111111010101001) && ({row_reg, col_reg}<18'b010111111010101011)) color_data = 12'b011111011110;
		if(({row_reg, col_reg}==18'b010111111010101011)) color_data = 12'b011011011110;
		if(({row_reg, col_reg}==18'b010111111010101100)) color_data = 12'b011111011110;
		if(({row_reg, col_reg}==18'b010111111010101101)) color_data = 12'b011011001110;
		if(({row_reg, col_reg}>=18'b010111111010101110) && ({row_reg, col_reg}<18'b010111111010110010)) color_data = 12'b011011011110;
		if(({row_reg, col_reg}==18'b010111111010110010)) color_data = 12'b011011001110;
		if(({row_reg, col_reg}==18'b010111111010110011)) color_data = 12'b010110111110;
		if(({row_reg, col_reg}==18'b010111111010110100)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}>=18'b010111111010110101) && ({row_reg, col_reg}<18'b010111111010110111)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b010111111010110111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b010111111010111000) && ({row_reg, col_reg}<18'b010111111010111010)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}>=18'b010111111010111010) && ({row_reg, col_reg}<18'b010111111010111101)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010111111010111101)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010111111010111110)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111111010111111)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b010111111011000000) && ({row_reg, col_reg}<18'b010111111011000010)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b010111111011000010)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b010111111011000011)) color_data = 12'b010010001110;
		if(({row_reg, col_reg}>=18'b010111111011000100) && ({row_reg, col_reg}<18'b010111111011000111)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}>=18'b010111111011000111) && ({row_reg, col_reg}<18'b010111111011001001)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010111111011001001)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b010111111011001010)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b010111111011001011)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010111111011001100)) color_data = 12'b010010001110;
		if(({row_reg, col_reg}==18'b010111111011001101)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}==18'b010111111011001110)) color_data = 12'b010010001110;
		if(({row_reg, col_reg}>=18'b010111111011001111) && ({row_reg, col_reg}<18'b010111111011011010)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}>=18'b010111111011011010) && ({row_reg, col_reg}<18'b010111111011011100)) color_data = 12'b010010001110;
		if(({row_reg, col_reg}>=18'b010111111011011100) && ({row_reg, col_reg}<18'b010111111011011110)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}==18'b010111111011011110)) color_data = 12'b010010011110;
		if(({row_reg, col_reg}>=18'b010111111011011111) && ({row_reg, col_reg}<18'b010111111011100010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010111111011100010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010111111011100011) && ({row_reg, col_reg}<18'b010111111011101001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b010111111011101001) && ({row_reg, col_reg}<18'b010111111011101011)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b010111111011101011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010111111011101100)) color_data = 12'b011010011110;
		if(({row_reg, col_reg}>=18'b010111111011101101) && ({row_reg, col_reg}<18'b010111111011110000)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010111111011110000)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b010111111011110001) && ({row_reg, col_reg}<18'b010111111011110011)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}>=18'b010111111011110011) && ({row_reg, col_reg}<18'b010111111011110110)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}==18'b010111111011110110)) color_data = 12'b010001111101;
		if(({row_reg, col_reg}>=18'b010111111011110111) && ({row_reg, col_reg}<18'b010111111011111010)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b010111111011111010)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b010111111011111011) && ({row_reg, col_reg}<18'b010111111011111101)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}>=18'b010111111011111101) && ({row_reg, col_reg}<18'b010111111011111111)) color_data = 12'b010010001110;
		if(({row_reg, col_reg}==18'b010111111011111111)) color_data = 12'b010110001110;
		if(({row_reg, col_reg}==18'b010111111100000000)) color_data = 12'b010110101110;
		if(({row_reg, col_reg}==18'b010111111100000001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010111111100000010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010111111100000011) && ({row_reg, col_reg}<18'b010111111100000110)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}==18'b010111111100000110)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}>=18'b010111111100000111) && ({row_reg, col_reg}<18'b010111111100001001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b010111111100001001)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b010111111100001010) && ({row_reg, col_reg}<18'b010111111100001100)) color_data = 12'b011010101110;

		if(({row_reg, col_reg}>=18'b010111111100001100) && ({row_reg, col_reg}<18'b011000000000000000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011000000000000000) && ({row_reg, col_reg}<18'b011000000000011000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011000000000011000)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==18'b011000000000011001)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011000000000011010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011000000000011011) && ({row_reg, col_reg}<18'b011000000000100000)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011000000000100000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011000000000100001) && ({row_reg, col_reg}<18'b011000000000100100)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011000000000100100)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==18'b011000000000100101)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}>=18'b011000000000100110) && ({row_reg, col_reg}<18'b011000000000101001)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011000000000101001)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000000000101010)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011000000000101011)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}==18'b011000000000101100)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000000000101101)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b011000000000101110)) color_data = 12'b010010011110;
		if(({row_reg, col_reg}==18'b011000000000101111)) color_data = 12'b010110101111;
		if(({row_reg, col_reg}>=18'b011000000000110000) && ({row_reg, col_reg}<18'b011000000000110010)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b011000000000110010) && ({row_reg, col_reg}<18'b011000000000111000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011000000000111000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b011000000000111001)) color_data = 12'b011110111110;
		if(({row_reg, col_reg}==18'b011000000000111010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b011000000000111011)) color_data = 12'b011110111110;
		if(({row_reg, col_reg}==18'b011000000000111100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011000000000111101)) color_data = 12'b011110111110;
		if(({row_reg, col_reg}>=18'b011000000000111110) && ({row_reg, col_reg}<18'b011000000001000000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011000000001000000)) color_data = 12'b010110101110;
		if(({row_reg, col_reg}==18'b011000000001000001)) color_data = 12'b001110011101;
		if(({row_reg, col_reg}==18'b011000000001000010)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b011000000001000011) && ({row_reg, col_reg}<18'b011000000001000101)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b011000000001000101)) color_data = 12'b001010011011;
		if(({row_reg, col_reg}==18'b011000000001000110)) color_data = 12'b011011011111;
		if(({row_reg, col_reg}==18'b011000000001000111)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b011000000001001000)) color_data = 12'b100011111110;
		if(({row_reg, col_reg}>=18'b011000000001001001) && ({row_reg, col_reg}<18'b011000000001001011)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b011000000001001011) && ({row_reg, col_reg}<18'b011000000001001101)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b011000000001001101) && ({row_reg, col_reg}<18'b011000000001001111)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b011000000001001111)) color_data = 12'b011011011110;
		if(({row_reg, col_reg}>=18'b011000000001010000) && ({row_reg, col_reg}<18'b011000000001010010)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b011000000001010010)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011000000001010011)) color_data = 12'b001010001101;
		if(({row_reg, col_reg}==18'b011000000001010100)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b011000000001010101)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b011000000001010110)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b011000000001010111)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b011000000001011000)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b011000000001011001) && ({row_reg, col_reg}<18'b011000000001011100)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b011000000001011100)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b011000000001011101)) color_data = 12'b001110011100;
		if(({row_reg, col_reg}==18'b011000000001011110)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}==18'b011000000001011111)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b011000000001100000)) color_data = 12'b100011111110;
		if(({row_reg, col_reg}>=18'b011000000001100001) && ({row_reg, col_reg}<18'b011000000001100100)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b011000000001100100)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}>=18'b011000000001100101) && ({row_reg, col_reg}<18'b011000000001100111)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b011000000001100111)) color_data = 12'b011110111110;
		if(({row_reg, col_reg}==18'b011000000001101000)) color_data = 12'b001101111010;
		if(({row_reg, col_reg}==18'b011000000001101001)) color_data = 12'b010001111010;
		if(({row_reg, col_reg}>=18'b011000000001101010) && ({row_reg, col_reg}<18'b011000000001101100)) color_data = 12'b001101111001;
		if(({row_reg, col_reg}==18'b011000000001101100)) color_data = 12'b011110111100;
		if(({row_reg, col_reg}==18'b011000000001101101)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}==18'b011000000001101110)) color_data = 12'b101011101111;
		if(({row_reg, col_reg}==18'b011000000001101111)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}==18'b011000000001110000)) color_data = 12'b100011101110;
		if(({row_reg, col_reg}==18'b011000000001110001)) color_data = 12'b010010011010;
		if(({row_reg, col_reg}==18'b011000000001110010)) color_data = 12'b001001111001;
		if(({row_reg, col_reg}==18'b011000000001110011)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b011000000001110100)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011000000001110101)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b011000000001110110)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011000000001110111) && ({row_reg, col_reg}<18'b011000000001111001)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011000000001111001)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011000000001111010)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}>=18'b011000000001111011) && ({row_reg, col_reg}<18'b011000000001111101)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b011000000001111101)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b011000000001111110) && ({row_reg, col_reg}<18'b011000000010000000)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b011000000010000000)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011000000010000001)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b011000000010000010)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b011000000010000011) && ({row_reg, col_reg}<18'b011000000010000111)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}>=18'b011000000010000111) && ({row_reg, col_reg}<18'b011000000010001001)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011000000010001001)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}>=18'b011000000010001010) && ({row_reg, col_reg}<18'b011000000010001101)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011000000010001101) && ({row_reg, col_reg}<18'b011000000010010000)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011000000010010000) && ({row_reg, col_reg}<18'b011000000010010011)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011000000010010011)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b011000000010010100) && ({row_reg, col_reg}<18'b011000000010011011)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011000000010011011) && ({row_reg, col_reg}<18'b011000000010011110)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}>=18'b011000000010011110) && ({row_reg, col_reg}<18'b011000000010100000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011000000010100000)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b011000000010100001) && ({row_reg, col_reg}<18'b011000000010100011)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b011000000010100011)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b011000000010100100)) color_data = 12'b001110001011;
		if(({row_reg, col_reg}==18'b011000000010100101)) color_data = 12'b010010011101;
		if(({row_reg, col_reg}==18'b011000000010100110)) color_data = 12'b010110101110;
		if(({row_reg, col_reg}==18'b011000000010100111)) color_data = 12'b010110101101;
		if(({row_reg, col_reg}==18'b011000000010101000)) color_data = 12'b010110101110;
		if(({row_reg, col_reg}==18'b011000000010101001)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==18'b011000000010101010)) color_data = 12'b010010011101;
		if(({row_reg, col_reg}>=18'b011000000010101011) && ({row_reg, col_reg}<18'b011000000010101111)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b011000000010101111)) color_data = 12'b001010001101;
		if(({row_reg, col_reg}==18'b011000000010110000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011000000010110001) && ({row_reg, col_reg}<18'b011000000010110011)) color_data = 12'b001010001101;
		if(({row_reg, col_reg}==18'b011000000010110011)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}>=18'b011000000010110100) && ({row_reg, col_reg}<18'b011000000010110110)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011000000010110110) && ({row_reg, col_reg}<18'b011000000010111000)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000000010111000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011000000010111001) && ({row_reg, col_reg}<18'b011000000010111011)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000000010111011)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b011000000010111100)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}==18'b011000000010111101)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b011000000010111110)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b011000000010111111)) color_data = 12'b001010001110;
		if(({row_reg, col_reg}==18'b011000000011000000)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011000000011000001)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b011000000011000010)) color_data = 12'b010110101111;
		if(({row_reg, col_reg}>=18'b011000000011000011) && ({row_reg, col_reg}<18'b011000000011000110)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011000000011000110)) color_data = 12'b010110011111;
		if(({row_reg, col_reg}==18'b011000000011000111)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}>=18'b011000000011001000) && ({row_reg, col_reg}<18'b011000000011001010)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000000011001010)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011000000011001011)) color_data = 12'b010010011110;
		if(({row_reg, col_reg}==18'b011000000011001100)) color_data = 12'b010110101111;
		if(({row_reg, col_reg}>=18'b011000000011001101) && ({row_reg, col_reg}<18'b011000000011001111)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b011000000011001111) && ({row_reg, col_reg}<18'b011000000011011111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011000000011011111)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==18'b011000000011100000)) color_data = 12'b011110101101;
		if(({row_reg, col_reg}>=18'b011000000011100001) && ({row_reg, col_reg}<18'b011000000011100011)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b011000000011100011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011000000011100100) && ({row_reg, col_reg}<18'b011000000011100110)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b011000000011100110) && ({row_reg, col_reg}<18'b011000000011101010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011000000011101010)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}>=18'b011000000011101011) && ({row_reg, col_reg}<18'b011000000011101101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011000000011101101)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}>=18'b011000000011101110) && ({row_reg, col_reg}<18'b011000000011110000)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b011000000011110000)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000000011110001)) color_data = 12'b010010001110;
		if(({row_reg, col_reg}==18'b011000000011110010)) color_data = 12'b010110101111;
		if(({row_reg, col_reg}>=18'b011000000011110011) && ({row_reg, col_reg}<18'b011000000011110110)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011000000011110110)) color_data = 12'b010010011110;
		if(({row_reg, col_reg}==18'b011000000011110111)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}>=18'b011000000011111000) && ({row_reg, col_reg}<18'b011000000011111011)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000000011111011)) color_data = 12'b010110101111;
		if(({row_reg, col_reg}>=18'b011000000011111100) && ({row_reg, col_reg}<18'b011000000100000000)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b011000000100000000) && ({row_reg, col_reg}<18'b011000000100000101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011000000100000101) && ({row_reg, col_reg}<18'b011000000100010000)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b011000000100010000) && ({row_reg, col_reg}<18'b011000001000011000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011000001000011000)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011000001000011001)) color_data = 12'b011110111111;
		if(({row_reg, col_reg}>=18'b011000001000011010) && ({row_reg, col_reg}<18'b011000001000100010)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b011000001000100010) && ({row_reg, col_reg}<18'b011000001000100100)) color_data = 12'b011010111111;
		if(({row_reg, col_reg}==18'b011000001000100100)) color_data = 12'b010110101111;
		if(({row_reg, col_reg}==18'b011000001000100101)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}==18'b011000001000100110)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000001000100111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011000001000101000)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}==18'b011000001000101001)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000001000101010)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011000001000101011)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000001000101100)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011000001000101101)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000001000101110)) color_data = 12'b010010011110;
		if(({row_reg, col_reg}==18'b011000001000101111)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011000001000110000)) color_data = 12'b011010111111;
		if(({row_reg, col_reg}==18'b011000001000110001)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b011000001000110010) && ({row_reg, col_reg}<18'b011000001000111010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011000001000111010) && ({row_reg, col_reg}<18'b011000001000111101)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}>=18'b011000001000111101) && ({row_reg, col_reg}<18'b011000001001000000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011000001001000000)) color_data = 12'b011010111111;
		if(({row_reg, col_reg}==18'b011000001001000001)) color_data = 12'b010010011110;
		if(({row_reg, col_reg}>=18'b011000001001000010) && ({row_reg, col_reg}<18'b011000001001000100)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011000001001000100)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b011000001001000101)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b011000001001000110)) color_data = 12'b011011011111;
		if(({row_reg, col_reg}==18'b011000001001000111)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b011000001001001000)) color_data = 12'b100011111110;
		if(({row_reg, col_reg}==18'b011000001001001001)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b011000001001001010) && ({row_reg, col_reg}<18'b011000001001001100)) color_data = 12'b100011111110;
		if(({row_reg, col_reg}==18'b011000001001001100)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b011000001001001101)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b011000001001001110)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b011000001001001111)) color_data = 12'b011111011110;
		if(({row_reg, col_reg}==18'b011000001001010000)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}>=18'b011000001001010001) && ({row_reg, col_reg}<18'b011000001001010101)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011000001001010101)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b011000001001010110)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b011000001001010111)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011000001001011000)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b011000001001011001)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b011000001001011010) && ({row_reg, col_reg}<18'b011000001001011100)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011000001001011100)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b011000001001011101)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b011000001001011110)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b011000001001011111)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b011000001001100000) && ({row_reg, col_reg}<18'b011000001001100100)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b011000001001100100)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}==18'b011000001001100101)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b011000001001100110)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b011000001001100111)) color_data = 12'b011111001110;
		if(({row_reg, col_reg}>=18'b011000001001101000) && ({row_reg, col_reg}<18'b011000001001101100)) color_data = 12'b001110001010;
		if(({row_reg, col_reg}==18'b011000001001101100)) color_data = 12'b011111001101;
		if(({row_reg, col_reg}==18'b011000001001101101)) color_data = 12'b101011111111;
		if(({row_reg, col_reg}==18'b011000001001101110)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b011000001001101111)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b011000001001110000)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b011000001001110001)) color_data = 12'b010010011011;
		if(({row_reg, col_reg}==18'b011000001001110010)) color_data = 12'b001010001010;
		if(({row_reg, col_reg}==18'b011000001001110011)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b011000001001110100)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b011000001001110101) && ({row_reg, col_reg}<18'b011000001001110111)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b011000001001110111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011000001001111000)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}>=18'b011000001001111001) && ({row_reg, col_reg}<18'b011000001001111100)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011000001001111100)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}>=18'b011000001001111101) && ({row_reg, col_reg}<18'b011000001001111111)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011000001001111111)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b011000001010000000)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b011000001010000001) && ({row_reg, col_reg}<18'b011000001010000011)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011000001010000011) && ({row_reg, col_reg}<18'b011000001010000110)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}>=18'b011000001010000110) && ({row_reg, col_reg}<18'b011000001010001100)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011000001010001100) && ({row_reg, col_reg}<18'b011000001010001111)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000001010001111)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b011000001010010000)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000001010010001)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b011000001010010010)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011000001010010011)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b011000001010010100)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011000001010010101)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b011000001010010110) && ({row_reg, col_reg}<18'b011000001010100000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011000001010100000) && ({row_reg, col_reg}<18'b011000001010100010)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b011000001010100010)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b011000001010100011)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b011000001010100100)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b011000001010100101)) color_data = 12'b010010011101;
		if(({row_reg, col_reg}>=18'b011000001010100110) && ({row_reg, col_reg}<18'b011000001010101000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011000001010101000)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==18'b011000001010101001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011000001010101010)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}>=18'b011000001010101011) && ({row_reg, col_reg}<18'b011000001010101111)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b011000001010101111) && ({row_reg, col_reg}<18'b011000001010110011)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011000001010110011)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011000001010110100) && ({row_reg, col_reg}<18'b011000001010110110)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011000001010110110) && ({row_reg, col_reg}<18'b011000001010111001)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000001010111001)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}>=18'b011000001010111010) && ({row_reg, col_reg}<18'b011000001010111100)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011000001010111100)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011000001010111101) && ({row_reg, col_reg}<18'b011000001010111111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011000001010111111)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b011000001011000000)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011000001011000001)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b011000001011000010)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b011000001011000011) && ({row_reg, col_reg}<18'b011000001011000110)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}==18'b011000001011000110)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==18'b011000001011000111)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}==18'b011000001011001000)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011000001011001001)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011000001011001010)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011000001011001011)) color_data = 12'b010010011110;
		if(({row_reg, col_reg}==18'b011000001011001100)) color_data = 12'b010110101111;
		if(({row_reg, col_reg}==18'b011000001011001101)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011000001011001110)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}>=18'b011000001011001111) && ({row_reg, col_reg}<18'b011000001011011001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011000001011011001)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}>=18'b011000001011011010) && ({row_reg, col_reg}<18'b011000001011100000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011000001011100000)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}>=18'b011000001011100001) && ({row_reg, col_reg}<18'b011000001011100100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011000001011100100)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b011000001011100101) && ({row_reg, col_reg}<18'b011000001011100111)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}==18'b011000001011100111)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011000001011101000) && ({row_reg, col_reg}<18'b011000001011101011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011000001011101011)) color_data = 12'b011110111110;
		if(({row_reg, col_reg}==18'b011000001011101100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011000001011101101)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}==18'b011000001011101110)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000001011101111)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b011000001011110000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011000001011110001)) color_data = 12'b010010011110;
		if(({row_reg, col_reg}>=18'b011000001011110010) && ({row_reg, col_reg}<18'b011000001011110100)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011000001011110100)) color_data = 12'b011010111111;
		if(({row_reg, col_reg}==18'b011000001011110101)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011000001011110110)) color_data = 12'b010010011110;
		if(({row_reg, col_reg}==18'b011000001011110111)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011000001011111000) && ({row_reg, col_reg}<18'b011000001011111010)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011000001011111010)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011000001011111011)) color_data = 12'b010110011111;
		if(({row_reg, col_reg}>=18'b011000001011111100) && ({row_reg, col_reg}<18'b011000001100000000)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b011000001100000000) && ({row_reg, col_reg}<18'b011000001100001000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011000001100001000) && ({row_reg, col_reg}<18'b011000001100010000)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b011000001100010000) && ({row_reg, col_reg}<18'b011000010000010011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011000010000010011)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011000010000010100) && ({row_reg, col_reg}<18'b011000010000010110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011000010000010110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011000010000010111) && ({row_reg, col_reg}<18'b011000010000011001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011000010000011001) && ({row_reg, col_reg}<18'b011000010000100011)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011000010000100011)) color_data = 12'b011010111111;
		if(({row_reg, col_reg}==18'b011000010000100100)) color_data = 12'b010110011111;
		if(({row_reg, col_reg}==18'b011000010000100101)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}>=18'b011000010000100110) && ({row_reg, col_reg}<18'b011000010000101000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011000010000101000)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000010000101001)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011000010000101010)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000010000101011)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b011000010000101100)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011000010000101101)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000010000101110)) color_data = 12'b010010011111;
		if(({row_reg, col_reg}==18'b011000010000101111)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011000010000110000)) color_data = 12'b011010111111;
		if(({row_reg, col_reg}>=18'b011000010000110001) && ({row_reg, col_reg}<18'b011000010000110011)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b011000010000110011) && ({row_reg, col_reg}<18'b011000010000110101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011000010000110101) && ({row_reg, col_reg}<18'b011000010000110111)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b011000010000110111) && ({row_reg, col_reg}<18'b011000010000111010)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}==18'b011000010000111010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011000010000111011)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011000010000111100) && ({row_reg, col_reg}<18'b011000010000111111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011000010000111111) && ({row_reg, col_reg}<18'b011000010001000001)) color_data = 12'b011010111111;
		if(({row_reg, col_reg}==18'b011000010001000001)) color_data = 12'b010010011110;
		if(({row_reg, col_reg}==18'b011000010001000010)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011000010001000011)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b011000010001000100)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b011000010001000101)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b011000010001000110)) color_data = 12'b011011001111;
		if(({row_reg, col_reg}==18'b011000010001000111)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b011000010001001000)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b011000010001001001) && ({row_reg, col_reg}<18'b011000010001001101)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b011000010001001101)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b011000010001001110)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b011000010001001111)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}==18'b011000010001010000)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b011000010001010001)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b011000010001010010)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}>=18'b011000010001010011) && ({row_reg, col_reg}<18'b011000010001011000)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b011000010001011000)) color_data = 12'b001010001101;
		if(({row_reg, col_reg}==18'b011000010001011001)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b011000010001011010)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011000010001011011)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b011000010001011100)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b011000010001011101)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b011000010001011110)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}>=18'b011000010001011111) && ({row_reg, col_reg}<18'b011000010001100100)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b011000010001100100)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b011000010001100101)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b011000010001100110)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b011000010001100111)) color_data = 12'b011011001110;
		if(({row_reg, col_reg}==18'b011000010001101000)) color_data = 12'b001010001010;
		if(({row_reg, col_reg}==18'b011000010001101001)) color_data = 12'b001110001010;
		if(({row_reg, col_reg}==18'b011000010001101010)) color_data = 12'b001010001010;
		if(({row_reg, col_reg}==18'b011000010001101011)) color_data = 12'b001010001001;
		if(({row_reg, col_reg}==18'b011000010001101100)) color_data = 12'b011011001101;
		if(({row_reg, col_reg}==18'b011000010001101101)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b011000010001101110)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b011000010001101111)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b011000010001110000)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b011000010001110001)) color_data = 12'b010010011100;
		if(({row_reg, col_reg}==18'b011000010001110010)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b011000010001110011)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b011000010001110100)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b011000010001110101) && ({row_reg, col_reg}<18'b011000010001111000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011000010001111000)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b011000010001111001)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011000010001111010)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b011000010001111011)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011000010001111100)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}>=18'b011000010001111101) && ({row_reg, col_reg}<18'b011000010001111111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011000010001111111)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}>=18'b011000010010000000) && ({row_reg, col_reg}<18'b011000010010000010)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011000010010000010)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}>=18'b011000010010000011) && ({row_reg, col_reg}<18'b011000010010000110)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011000010010000110)) color_data = 12'b001010001101;
		if(({row_reg, col_reg}>=18'b011000010010000111) && ({row_reg, col_reg}<18'b011000010010001001)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b011000010010001001) && ({row_reg, col_reg}<18'b011000010010001011)) color_data = 12'b001010001101;
		if(({row_reg, col_reg}>=18'b011000010010001011) && ({row_reg, col_reg}<18'b011000010010001101)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011000010010001101)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011000010010001110) && ({row_reg, col_reg}<18'b011000010010010000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011000010010010000)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b011000010010010001)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b011000010010010010)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b011000010010010011)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b011000010010010100)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b011000010010010101)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b011000010010010110) && ({row_reg, col_reg}<18'b011000010010011101)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011000010010011101) && ({row_reg, col_reg}<18'b011000010010100001)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000010010100001)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011000010010100010) && ({row_reg, col_reg}<18'b011000010010100100)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000010010100100)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b011000010010100101)) color_data = 12'b010010011110;
		if(({row_reg, col_reg}>=18'b011000010010100110) && ({row_reg, col_reg}<18'b011000010010101000)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011000010010101000)) color_data = 12'b011010111111;
		if(({row_reg, col_reg}==18'b011000010010101001)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011000010010101010)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}==18'b011000010010101011)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}>=18'b011000010010101100) && ({row_reg, col_reg}<18'b011000010010101110)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000010010101110)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}>=18'b011000010010101111) && ({row_reg, col_reg}<18'b011000010010110001)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011000010010110001) && ({row_reg, col_reg}<18'b011000010010111011)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000010010111011)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b011000010010111100) && ({row_reg, col_reg}<18'b011000010010111110)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b011000010010111110)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000010010111111)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b011000010011000000)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011000010011000001)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b011000010011000010)) color_data = 12'b010110101110;
		if(({row_reg, col_reg}>=18'b011000010011000011) && ({row_reg, col_reg}<18'b011000010011000110)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011000010011000110)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==18'b011000010011000111)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b011000010011001000)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b011000010011001001) && ({row_reg, col_reg}<18'b011000010011001011)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b011000010011001011)) color_data = 12'b010010011101;
		if(({row_reg, col_reg}==18'b011000010011001100)) color_data = 12'b010110101110;
		if(({row_reg, col_reg}==18'b011000010011001101)) color_data = 12'b011110111111;
		if(({row_reg, col_reg}==18'b011000010011001110)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}>=18'b011000010011001111) && ({row_reg, col_reg}<18'b011000010011100000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011000010011100000) && ({row_reg, col_reg}<18'b011000010011100011)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011000010011100011) && ({row_reg, col_reg}<18'b011000010011101011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011000010011101011)) color_data = 12'b011110111111;
		if(({row_reg, col_reg}==18'b011000010011101100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011000010011101101)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}>=18'b011000010011101110) && ({row_reg, col_reg}<18'b011000010011110000)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000010011110000)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011000010011110001)) color_data = 12'b010010011110;
		if(({row_reg, col_reg}>=18'b011000010011110010) && ({row_reg, col_reg}<18'b011000010011110110)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011000010011110110)) color_data = 12'b010010011101;
		if(({row_reg, col_reg}>=18'b011000010011110111) && ({row_reg, col_reg}<18'b011000010011111001)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}>=18'b011000010011111001) && ({row_reg, col_reg}<18'b011000010011111011)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000010011111011)) color_data = 12'b010110101110;
		if(({row_reg, col_reg}>=18'b011000010011111100) && ({row_reg, col_reg}<18'b011000010011111111)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b011000010011111111) && ({row_reg, col_reg}<18'b011000010100000101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011000010100000101) && ({row_reg, col_reg}<18'b011000010100010000)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b011000010100010000) && ({row_reg, col_reg}<18'b011000011000010011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011000011000010011)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011000011000010100) && ({row_reg, col_reg}<18'b011000011000011010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011000011000011010) && ({row_reg, col_reg}<18'b011000011000100100)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011000011000100100)) color_data = 12'b010110101111;
		if(({row_reg, col_reg}==18'b011000011000100101)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}==18'b011000011000100110)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011000011000100111) && ({row_reg, col_reg}<18'b011000011000101001)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000011000101001)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011000011000101010)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}==18'b011000011000101011)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000011000101100)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011000011000101101)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000011000101110)) color_data = 12'b010010011111;
		if(({row_reg, col_reg}==18'b011000011000101111)) color_data = 12'b010110101111;
		if(({row_reg, col_reg}>=18'b011000011000110000) && ({row_reg, col_reg}<18'b011000011000110111)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011000011000110111)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}>=18'b011000011000111000) && ({row_reg, col_reg}<18'b011000011000111011)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011000011000111011)) color_data = 12'b011110111111;
		if(({row_reg, col_reg}>=18'b011000011000111100) && ({row_reg, col_reg}<18'b011000011001000000)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011000011001000000)) color_data = 12'b010110101111;
		if(({row_reg, col_reg}==18'b011000011001000001)) color_data = 12'b010010001110;
		if(({row_reg, col_reg}>=18'b011000011001000010) && ({row_reg, col_reg}<18'b011000011001000100)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000011001000100)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011000011001000101)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b011000011001000110)) color_data = 12'b011111001111;
		if(({row_reg, col_reg}>=18'b011000011001000111) && ({row_reg, col_reg}<18'b011000011001001101)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b011000011001001101)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b011000011001001110)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b011000011001001111)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}>=18'b011000011001010000) && ({row_reg, col_reg}<18'b011000011001010101)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b011000011001010101)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}>=18'b011000011001010110) && ({row_reg, col_reg}<18'b011000011001011000)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}>=18'b011000011001011000) && ({row_reg, col_reg}<18'b011000011001011010)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b011000011001011010)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011000011001011011)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b011000011001011100)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b011000011001011101)) color_data = 12'b001110011100;
		if(({row_reg, col_reg}==18'b011000011001011110)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b011000011001011111)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b011000011001100000) && ({row_reg, col_reg}<18'b011000011001100011)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b011000011001100011) && ({row_reg, col_reg}<18'b011000011001100101)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b011000011001100101) && ({row_reg, col_reg}<18'b011000011001100111)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b011000011001100111)) color_data = 12'b011011011110;
		if(({row_reg, col_reg}>=18'b011000011001101000) && ({row_reg, col_reg}<18'b011000011001101010)) color_data = 12'b001010001010;
		if(({row_reg, col_reg}>=18'b011000011001101010) && ({row_reg, col_reg}<18'b011000011001101100)) color_data = 12'b001010011010;
		if(({row_reg, col_reg}==18'b011000011001101100)) color_data = 12'b010111001101;
		if(({row_reg, col_reg}>=18'b011000011001101101) && ({row_reg, col_reg}<18'b011000011001110000)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b011000011001110000)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b011000011001110001)) color_data = 12'b010010101100;
		if(({row_reg, col_reg}==18'b011000011001110010)) color_data = 12'b001001111010;
		if(({row_reg, col_reg}==18'b011000011001110011)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}>=18'b011000011001110100) && ({row_reg, col_reg}<18'b011000011001110111)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011000011001110111)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}>=18'b011000011001111000) && ({row_reg, col_reg}<18'b011000011001111010)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b011000011001111010)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011000011001111011)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011000011001111100)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b011000011001111101) && ({row_reg, col_reg}<18'b011000011001111111)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b011000011001111111)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b011000011010000000)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}>=18'b011000011010000001) && ({row_reg, col_reg}<18'b011000011010000011)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011000011010000011)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b011000011010000100) && ({row_reg, col_reg}<18'b011000011010000111)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}>=18'b011000011010000111) && ({row_reg, col_reg}<18'b011000011010001001)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b011000011010001001)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b011000011010001010)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b011000011010001011)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b011000011010001100)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b011000011010001101)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b011000011010001110)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011000011010001111)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}==18'b011000011010010000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011000011010010001)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b011000011010010010) && ({row_reg, col_reg}<18'b011000011010010100)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}>=18'b011000011010010100) && ({row_reg, col_reg}<18'b011000011010011100)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011000011010011100)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000011010011101)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b011000011010011110)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000011010011111)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}>=18'b011000011010100000) && ({row_reg, col_reg}<18'b011000011010100011)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011000011010100011) && ({row_reg, col_reg}<18'b011000011010100101)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b011000011010100101)) color_data = 12'b010110001110;
		if(({row_reg, col_reg}==18'b011000011010100110)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011000011010100111)) color_data = 12'b011110111111;
		if(({row_reg, col_reg}==18'b011000011010101000)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}==18'b011000011010101001)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011000011010101010)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}>=18'b011000011010101011) && ({row_reg, col_reg}<18'b011000011010111000)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000011010111000)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b011000011010111001)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011000011010111010) && ({row_reg, col_reg}<18'b011000011011000001)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b011000011011000001)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}==18'b011000011011000010)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==18'b011000011011000011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011000011011000100) && ({row_reg, col_reg}<18'b011000011011000110)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011000011011000110)) color_data = 12'b011010011110;
		if(({row_reg, col_reg}==18'b011000011011000111)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}>=18'b011000011011001000) && ({row_reg, col_reg}<18'b011000011011001010)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b011000011011001010)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b011000011011001011)) color_data = 12'b010010011110;
		if(({row_reg, col_reg}==18'b011000011011001100)) color_data = 12'b010110101110;
		if(({row_reg, col_reg}==18'b011000011011001101)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b011000011011001110) && ({row_reg, col_reg}<18'b011000011011100110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011000011011100110) && ({row_reg, col_reg}<18'b011000011011101000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011000011011101000) && ({row_reg, col_reg}<18'b011000011011101100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011000011011101100)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==18'b011000011011101101)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}>=18'b011000011011101110) && ({row_reg, col_reg}<18'b011000011011110000)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b011000011011110000)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000011011110001)) color_data = 12'b010010011110;
		if(({row_reg, col_reg}>=18'b011000011011110010) && ({row_reg, col_reg}<18'b011000011011110101)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011000011011110101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011000011011110110)) color_data = 12'b010110011101;
		if(({row_reg, col_reg}==18'b011000011011110111)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}>=18'b011000011011111000) && ({row_reg, col_reg}<18'b011000011011111011)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}>=18'b011000011011111011) && ({row_reg, col_reg}<18'b011000011011111101)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b011000011011111101) && ({row_reg, col_reg}<18'b011000011011111111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011000011011111111)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}>=18'b011000011100000000) && ({row_reg, col_reg}<18'b011000011100000110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011000011100000110) && ({row_reg, col_reg}<18'b011000011100001110)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b011000011100001110) && ({row_reg, col_reg}<18'b011000100000010000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011000100000010000) && ({row_reg, col_reg}<18'b011000100000010100)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011000100000010100) && ({row_reg, col_reg}<18'b011000100000010110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011000100000010110) && ({row_reg, col_reg}<18'b011000100000011000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b011000100000011000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011000100000011001) && ({row_reg, col_reg}<18'b011000100000011011)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011000100000011011)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}>=18'b011000100000011100) && ({row_reg, col_reg}<18'b011000100000100001)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}==18'b011000100000100001)) color_data = 12'b010010001110;
		if(({row_reg, col_reg}==18'b011000100000100010)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b011000100000100011)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}==18'b011000100000100100)) color_data = 12'b010010001110;
		if(({row_reg, col_reg}>=18'b011000100000100101) && ({row_reg, col_reg}<18'b011000100000100111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011000100000100111)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b011000100000101000)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011000100000101001) && ({row_reg, col_reg}<18'b011000100000101011)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011000100000101011)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000100000101100)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011000100000101101)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000100000101110)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}>=18'b011000100000101111) && ({row_reg, col_reg}<18'b011000100000110001)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}>=18'b011000100000110001) && ({row_reg, col_reg}<18'b011000100000110011)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}>=18'b011000100000110011) && ({row_reg, col_reg}<18'b011000100000111111)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}>=18'b011000100000111111) && ({row_reg, col_reg}<18'b011000100001000001)) color_data = 12'b010010001110;
		if(({row_reg, col_reg}==18'b011000100001000001)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b011000100001000010) && ({row_reg, col_reg}<18'b011000100001000100)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000100001000100)) color_data = 12'b001001101100;
		if(({row_reg, col_reg}==18'b011000100001000101)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011000100001000110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011000100001000111)) color_data = 12'b011111001111;
		if(({row_reg, col_reg}>=18'b011000100001001000) && ({row_reg, col_reg}<18'b011000100001001100)) color_data = 12'b011011001101;
		if(({row_reg, col_reg}==18'b011000100001001100)) color_data = 12'b011111001101;
		if(({row_reg, col_reg}>=18'b011000100001001101) && ({row_reg, col_reg}<18'b011000100001010000)) color_data = 12'b011111001110;
		if(({row_reg, col_reg}==18'b011000100001010000)) color_data = 12'b011011001110;
		if(({row_reg, col_reg}==18'b011000100001010001)) color_data = 12'b011111011110;
		if(({row_reg, col_reg}>=18'b011000100001010010) && ({row_reg, col_reg}<18'b011000100001011100)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}==18'b011000100001011100)) color_data = 12'b011111011110;
		if(({row_reg, col_reg}==18'b011000100001011101)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}==18'b011000100001011110)) color_data = 12'b010110111101;
		if(({row_reg, col_reg}==18'b011000100001011111)) color_data = 12'b010010101100;
		if(({row_reg, col_reg}==18'b011000100001100000)) color_data = 12'b010010101101;
		if(({row_reg, col_reg}==18'b011000100001100001)) color_data = 12'b010010101100;
		if(({row_reg, col_reg}==18'b011000100001100010)) color_data = 12'b010110111100;
		if(({row_reg, col_reg}==18'b011000100001100011)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b011000100001100100)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b011000100001100101)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b011000100001100110)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b011000100001100111)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b011000100001101000)) color_data = 12'b011011001101;
		if(({row_reg, col_reg}>=18'b011000100001101001) && ({row_reg, col_reg}<18'b011000100001101100)) color_data = 12'b011011011110;
		if(({row_reg, col_reg}>=18'b011000100001101100) && ({row_reg, col_reg}<18'b011000100001101110)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b011000100001101110)) color_data = 12'b011111111111;
		if(({row_reg, col_reg}>=18'b011000100001101111) && ({row_reg, col_reg}<18'b011000100001110001)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b011000100001110001)) color_data = 12'b011111101111;
		if(({row_reg, col_reg}==18'b011000100001110010)) color_data = 12'b011011011110;
		if(({row_reg, col_reg}==18'b011000100001110011)) color_data = 12'b011011011111;
		if(({row_reg, col_reg}>=18'b011000100001110100) && ({row_reg, col_reg}<18'b011000100001110110)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}==18'b011000100001110110)) color_data = 12'b100011011111;
		if(({row_reg, col_reg}==18'b011000100001110111)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}>=18'b011000100001111000) && ({row_reg, col_reg}<18'b011000100001111010)) color_data = 12'b011111001111;
		if(({row_reg, col_reg}==18'b011000100001111010)) color_data = 12'b010110101110;
		if(({row_reg, col_reg}==18'b011000100001111011)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011000100001111100)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}>=18'b011000100001111101) && ({row_reg, col_reg}<18'b011000100010000001)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b011000100010000001)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011000100010000010)) color_data = 12'b001010001101;
		if(({row_reg, col_reg}==18'b011000100010000011)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b011000100010000100)) color_data = 12'b010110111110;
		if(({row_reg, col_reg}==18'b011000100010000101)) color_data = 12'b011011001111;
		if(({row_reg, col_reg}>=18'b011000100010000110) && ({row_reg, col_reg}<18'b011000100010001100)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}==18'b011000100010001100)) color_data = 12'b011111001111;
		if(({row_reg, col_reg}==18'b011000100010001101)) color_data = 12'b011010111111;
		if(({row_reg, col_reg}==18'b011000100010001110)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b011000100010001111)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011000100010010000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011000100010010001)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b011000100010010010) && ({row_reg, col_reg}<18'b011000100010010100)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}>=18'b011000100010010100) && ({row_reg, col_reg}<18'b011000100010010111)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b011000100010010111) && ({row_reg, col_reg}<18'b011000100010011011)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000100010011011)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b011000100010011100)) color_data = 12'b010010011110;
		if(({row_reg, col_reg}==18'b011000100010011101)) color_data = 12'b010110011111;
		if(({row_reg, col_reg}==18'b011000100010011110)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==18'b011000100010011111)) color_data = 12'b010110011111;
		if(({row_reg, col_reg}>=18'b011000100010100000) && ({row_reg, col_reg}<18'b011000100010100100)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}>=18'b011000100010100100) && ({row_reg, col_reg}<18'b011000100010100110)) color_data = 12'b011010011110;
		if(({row_reg, col_reg}==18'b011000100010100110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011000100010100111) && ({row_reg, col_reg}<18'b011000100010101001)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}==18'b011000100010101001)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011000100010101010)) color_data = 12'b011010011110;
		if(({row_reg, col_reg}>=18'b011000100010101011) && ({row_reg, col_reg}<18'b011000100010101110)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}>=18'b011000100010101110) && ({row_reg, col_reg}<18'b011000100010110011)) color_data = 12'b010110011111;
		if(({row_reg, col_reg}==18'b011000100010110011)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==18'b011000100010110100)) color_data = 12'b010110011111;
		if(({row_reg, col_reg}>=18'b011000100010110101) && ({row_reg, col_reg}<18'b011000100011000000)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==18'b011000100011000000)) color_data = 12'b010110011101;
		if(({row_reg, col_reg}==18'b011000100011000001)) color_data = 12'b010110101110;
		if(({row_reg, col_reg}>=18'b011000100011000010) && ({row_reg, col_reg}<18'b011000100011000100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011000100011000100) && ({row_reg, col_reg}<18'b011000100011000110)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}==18'b011000100011000110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011000100011000111) && ({row_reg, col_reg}<18'b011000100011001011)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==18'b011000100011001011)) color_data = 12'b010110101110;
		if(({row_reg, col_reg}==18'b011000100011001100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011000100011001101)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b011000100011001110) && ({row_reg, col_reg}<18'b011000100011011000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011000100011011000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011000100011011001) && ({row_reg, col_reg}<18'b011000100011101011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011000100011101011)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}==18'b011000100011101100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011000100011101101) && ({row_reg, col_reg}<18'b011000100011110010)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}>=18'b011000100011110010) && ({row_reg, col_reg}<18'b011000100011110101)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b011000100011110101) && ({row_reg, col_reg}<18'b011000100011110111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011000100011110111) && ({row_reg, col_reg}<18'b011000100011111011)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==18'b011000100011111011)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b011000100011111100) && ({row_reg, col_reg}<18'b011000100011111111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011000100011111111) && ({row_reg, col_reg}<18'b011000100100000011)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011000100100000011) && ({row_reg, col_reg}<18'b011000100100000111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011000100100000111) && ({row_reg, col_reg}<18'b011000100100001011)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b011000100100001011) && ({row_reg, col_reg}<18'b011000101000010000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011000101000010000) && ({row_reg, col_reg}<18'b011000101000010101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011000101000010101) && ({row_reg, col_reg}<18'b011000101000011001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011000101000011001) && ({row_reg, col_reg}<18'b011000101000011011)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011000101000011011)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}>=18'b011000101000011100) && ({row_reg, col_reg}<18'b011000101000011110)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b011000101000011110)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000101000011111)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}>=18'b011000101000100000) && ({row_reg, col_reg}<18'b011000101000100010)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000101000100010)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011000101000100011)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011000101000100100)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011000101000100101) && ({row_reg, col_reg}<18'b011000101000100111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011000101000100111)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}==18'b011000101000101000)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000101000101001)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011000101000101010) && ({row_reg, col_reg}<18'b011000101000101100)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011000101000101100) && ({row_reg, col_reg}<18'b011000101000110011)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011000101000110011) && ({row_reg, col_reg}<18'b011000101000110101)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}>=18'b011000101000110101) && ({row_reg, col_reg}<18'b011000101000111010)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011000101000111010) && ({row_reg, col_reg}<18'b011000101000111101)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}>=18'b011000101000111101) && ({row_reg, col_reg}<18'b011000101000111111)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000101000111111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011000101001000000) && ({row_reg, col_reg}<18'b011000101001000011)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000101001000011)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b011000101001000100)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000101001000101)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b011000101001000110)) color_data = 12'b010110101110;
		if(({row_reg, col_reg}==18'b011000101001000111)) color_data = 12'b011010111111;
		if(({row_reg, col_reg}==18'b011000101001001000)) color_data = 12'b010110101101;
		if(({row_reg, col_reg}>=18'b011000101001001001) && ({row_reg, col_reg}<18'b011000101001001011)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}==18'b011000101001001011)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}==18'b011000101001001100)) color_data = 12'b010110101101;
		if(({row_reg, col_reg}==18'b011000101001001101)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}==18'b011000101001001110)) color_data = 12'b010110101100;
		if(({row_reg, col_reg}==18'b011000101001001111)) color_data = 12'b011111001110;
		if(({row_reg, col_reg}>=18'b011000101001010000) && ({row_reg, col_reg}<18'b011000101001010100)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b011000101001010100) && ({row_reg, col_reg}<18'b011000101001010110)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b011000101001010110) && ({row_reg, col_reg}<18'b011000101001011101)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b011000101001011101)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b011000101001011110)) color_data = 12'b001110011011;
		if(({row_reg, col_reg}==18'b011000101001011111)) color_data = 12'b001001111010;
		if(({row_reg, col_reg}==18'b011000101001100000)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b011000101001100001)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b011000101001100010)) color_data = 12'b001110011011;
		if(({row_reg, col_reg}==18'b011000101001100011)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b011000101001100100) && ({row_reg, col_reg}<18'b011000101001100111)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b011000101001100111) && ({row_reg, col_reg}<18'b011000101001110001)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b011000101001110001)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b011000101001110010)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b011000101001110011)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b011000101001110100)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b011000101001110101)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}>=18'b011000101001110110) && ({row_reg, col_reg}<18'b011000101001111010)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b011000101001111010)) color_data = 12'b011111001111;
		if(({row_reg, col_reg}==18'b011000101001111011)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}>=18'b011000101001111100) && ({row_reg, col_reg}<18'b011000101010000000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011000101010000000)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b011000101010000001)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}==18'b011000101010000010)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b011000101010000011)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b011000101010000100)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}>=18'b011000101010000101) && ({row_reg, col_reg}<18'b011000101010001101)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b011000101010001101)) color_data = 12'b011111001111;
		if(({row_reg, col_reg}==18'b011000101010001110)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b011000101010001111)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011000101010010000)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b011000101010010001)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}>=18'b011000101010010010) && ({row_reg, col_reg}<18'b011000101010011000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011000101010011000) && ({row_reg, col_reg}<18'b011000101010011011)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000101010011011)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b011000101010011100)) color_data = 12'b010110101111;
		if(({row_reg, col_reg}==18'b011000101010011101)) color_data = 12'b011010111111;
		if(({row_reg, col_reg}>=18'b011000101010011110) && ({row_reg, col_reg}<18'b011000101010100010)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011000101010100010)) color_data = 12'b011110111111;
		if(({row_reg, col_reg}>=18'b011000101010100011) && ({row_reg, col_reg}<18'b011000101010100101)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}==18'b011000101010100101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011000101010100110) && ({row_reg, col_reg}<18'b011000101010101001)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b011000101010101001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011000101010101010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b011000101010101011)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}>=18'b011000101010101100) && ({row_reg, col_reg}<18'b011000101010111110)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011000101010111110)) color_data = 12'b011010111111;
		if(({row_reg, col_reg}==18'b011000101010111111)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b011000101011000000) && ({row_reg, col_reg}<18'b011000101011000010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011000101011000010)) color_data = 12'b011110111111;
		if(({row_reg, col_reg}>=18'b011000101011000011) && ({row_reg, col_reg}<18'b011000101011001000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011000101011001000) && ({row_reg, col_reg}<18'b011000101011001101)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011000101011001101)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}==18'b011000101011001110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011000101011001111) && ({row_reg, col_reg}<18'b011000101011101011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011000101011101011)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011000101011101100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011000101011101101)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b011000101011101110) && ({row_reg, col_reg}<18'b011000101011110000)) color_data = 12'b011110111111;
		if(({row_reg, col_reg}>=18'b011000101011110000) && ({row_reg, col_reg}<18'b011000101011110011)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b011000101011110011) && ({row_reg, col_reg}<18'b011000101011110110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011000101011110110) && ({row_reg, col_reg}<18'b011000101011111001)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b011000101011111001) && ({row_reg, col_reg}<18'b011000101011111011)) color_data = 12'b011110111111;
		if(({row_reg, col_reg}>=18'b011000101011111011) && ({row_reg, col_reg}<18'b011000101011111110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011000101011111110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011000101011111111) && ({row_reg, col_reg}<18'b011000101100000101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011000101100000101) && ({row_reg, col_reg}<18'b011000101100001000)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b011000101100001000) && ({row_reg, col_reg}<18'b011000110000010000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011000110000010000) && ({row_reg, col_reg}<18'b011000110000010101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011000110000010101) && ({row_reg, col_reg}<18'b011000110000011000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011000110000011000) && ({row_reg, col_reg}<18'b011000110000011011)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011000110000011011)) color_data = 12'b010010001110;
		if(({row_reg, col_reg}==18'b011000110000011100)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000110000011101)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b011000110000011110) && ({row_reg, col_reg}<18'b011000110000100100)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000110000100100)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}>=18'b011000110000100101) && ({row_reg, col_reg}<18'b011000110000100111)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000110000100111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011000110000101000) && ({row_reg, col_reg}<18'b011000110000101010)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000110000101010)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}>=18'b011000110000101011) && ({row_reg, col_reg}<18'b011000110000101110)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011000110000101110)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b011000110000101111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011000110000110000) && ({row_reg, col_reg}<18'b011000110000110010)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000110000110010)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}>=18'b011000110000110011) && ({row_reg, col_reg}<18'b011000110000111111)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000110000111111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011000110001000000)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011000110001000001) && ({row_reg, col_reg}<18'b011000110001000011)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b011000110001000011) && ({row_reg, col_reg}<18'b011000110001000110)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000110001000110)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==18'b011000110001000111)) color_data = 12'b011010111111;
		if(({row_reg, col_reg}==18'b011000110001001000)) color_data = 12'b010110101110;
		if(({row_reg, col_reg}>=18'b011000110001001001) && ({row_reg, col_reg}<18'b011000110001001100)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==18'b011000110001001100)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}==18'b011000110001001101)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==18'b011000110001001110)) color_data = 12'b010110101100;
		if(({row_reg, col_reg}==18'b011000110001001111)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==18'b011000110001010000)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b011000110001010001)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b011000110001010010)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}>=18'b011000110001010011) && ({row_reg, col_reg}<18'b011000110001010110)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b011000110001010110)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b011000110001010111) && ({row_reg, col_reg}<18'b011000110001011010)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b011000110001011010)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b011000110001011011)) color_data = 12'b100011101110;
		if(({row_reg, col_reg}==18'b011000110001011100)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b011000110001011101)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b011000110001011110)) color_data = 12'b001110001011;
		if(({row_reg, col_reg}==18'b011000110001011111)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b011000110001100000)) color_data = 12'b001010001101;
		if(({row_reg, col_reg}==18'b011000110001100001)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011000110001100010)) color_data = 12'b010010101100;
		if(({row_reg, col_reg}==18'b011000110001100011)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b011000110001100100)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b011000110001100101) && ({row_reg, col_reg}<18'b011000110001100111)) color_data = 12'b100011111110;
		if(({row_reg, col_reg}>=18'b011000110001100111) && ({row_reg, col_reg}<18'b011000110001101001)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b011000110001101001)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b011000110001101010) && ({row_reg, col_reg}<18'b011000110001110001)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b011000110001110001)) color_data = 12'b100011111110;
		if(({row_reg, col_reg}>=18'b011000110001110010) && ({row_reg, col_reg}<18'b011000110001110101)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b011000110001110101)) color_data = 12'b100011111110;
		if(({row_reg, col_reg}>=18'b011000110001110110) && ({row_reg, col_reg}<18'b011000110001111000)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b011000110001111000)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b011000110001111001)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b011000110001111010)) color_data = 12'b011011001110;
		if(({row_reg, col_reg}==18'b011000110001111011)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b011000110001111100)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b011000110001111101)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}>=18'b011000110001111110) && ({row_reg, col_reg}<18'b011000110010000001)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011000110010000001)) color_data = 12'b001010001101;
		if(({row_reg, col_reg}==18'b011000110010000010)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011000110010000011)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b011000110010000100)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}==18'b011000110010000101)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b011000110010000110)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b011000110010000111)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b011000110010001000)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b011000110010001001)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b011000110010001010)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b011000110010001011)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b011000110010001100)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b011000110010001101)) color_data = 12'b011111001111;
		if(({row_reg, col_reg}==18'b011000110010001110)) color_data = 12'b001110001011;
		if(({row_reg, col_reg}==18'b011000110010001111)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011000110010010000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011000110010010001)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000110010010010)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011000110010010011)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000110010010100)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011000110010010101) && ({row_reg, col_reg}<18'b011000110010011010)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011000110010011010) && ({row_reg, col_reg}<18'b011000110010011100)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b011000110010011100)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==18'b011000110010011101)) color_data = 12'b011010111111;
		if(({row_reg, col_reg}>=18'b011000110010011110) && ({row_reg, col_reg}<18'b011000110010100011)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b011000110010100011) && ({row_reg, col_reg}<18'b011000110010101111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011000110010101111)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b011000110010110000) && ({row_reg, col_reg}<18'b011000110011001001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011000110011001001) && ({row_reg, col_reg}<18'b011000110011001011)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011000110011001011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011000110011001100)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011000110011001101) && ({row_reg, col_reg}<18'b011000110011001111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011000110011001111)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011000110011010000) && ({row_reg, col_reg}<18'b011000110011111000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011000110011111000)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b011000110011111001) && ({row_reg, col_reg}<18'b011000110011111100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011000110011111100)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b011000110011111101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011000110011111110) && ({row_reg, col_reg}<18'b011000110100000000)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b011000110100000000) && ({row_reg, col_reg}<18'b011000111000010000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011000111000010000) && ({row_reg, col_reg}<18'b011000111000010010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b011000111000010010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011000111000010011)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011000111000010100) && ({row_reg, col_reg}<18'b011000111000010110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011000111000010110) && ({row_reg, col_reg}<18'b011000111000011000)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011000111000011000)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}==18'b011000111000011001)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011000111000011010)) color_data = 12'b011110111111;
		if(({row_reg, col_reg}==18'b011000111000011011)) color_data = 12'b010010001110;
		if(({row_reg, col_reg}>=18'b011000111000011100) && ({row_reg, col_reg}<18'b011000111000100000)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000111000100000)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b011000111000100001)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}==18'b011000111000100010)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000111000100011)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011000111000100100) && ({row_reg, col_reg}<18'b011000111000100110)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011000111000100110) && ({row_reg, col_reg}<18'b011000111000101100)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011000111000101100)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000111000101101)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011000111000101110)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b011000111000101111) && ({row_reg, col_reg}<18'b011000111000110001)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011000111000110001) && ({row_reg, col_reg}<18'b011000111001000011)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000111001000011)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011000111001000100)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000111001000101)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011000111001000110)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==18'b011000111001000111)) color_data = 12'b011010111111;
		if(({row_reg, col_reg}==18'b011000111001001000)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b011000111001001001) && ({row_reg, col_reg}<18'b011000111001001100)) color_data = 12'b011010111111;
		if(({row_reg, col_reg}==18'b011000111001001100)) color_data = 12'b010110101110;
		if(({row_reg, col_reg}==18'b011000111001001101)) color_data = 12'b011011001111;
		if(({row_reg, col_reg}==18'b011000111001001110)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==18'b011000111001001111)) color_data = 12'b011111001111;
		if(({row_reg, col_reg}>=18'b011000111001010000) && ({row_reg, col_reg}<18'b011000111001010011)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b011000111001010011) && ({row_reg, col_reg}<18'b011000111001010101)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b011000111001010101)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b011000111001010110)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b011000111001010111) && ({row_reg, col_reg}<18'b011000111001011101)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b011000111001011101)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b011000111001011110)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b011000111001011111)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011000111001100000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011000111001100001)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011000111001100010)) color_data = 12'b010010101101;
		if(({row_reg, col_reg}>=18'b011000111001100011) && ({row_reg, col_reg}<18'b011000111001101001)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b011000111001101001) && ({row_reg, col_reg}<18'b011000111001110000)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b011000111001110000) && ({row_reg, col_reg}<18'b011000111001110010)) color_data = 12'b100011111110;
		if(({row_reg, col_reg}>=18'b011000111001110010) && ({row_reg, col_reg}<18'b011000111001110100)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b011000111001110100) && ({row_reg, col_reg}<18'b011000111001111010)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b011000111001111010)) color_data = 12'b011111001111;
		if(({row_reg, col_reg}==18'b011000111001111011)) color_data = 12'b001001111010;
		if(({row_reg, col_reg}==18'b011000111001111100)) color_data = 12'b000101111010;
		if(({row_reg, col_reg}==18'b011000111001111101)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b011000111001111110)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b011000111001111111)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011000111010000000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011000111010000001)) color_data = 12'b001010001101;
		if(({row_reg, col_reg}==18'b011000111010000010)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011000111010000011)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b011000111010000100)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}>=18'b011000111010000101) && ({row_reg, col_reg}<18'b011000111010001101)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b011000111010001101)) color_data = 12'b011111001111;
		if(({row_reg, col_reg}==18'b011000111010001110)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b011000111010001111)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b011000111010010000) && ({row_reg, col_reg}<18'b011000111010010010)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011000111010010010)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011000111010010011) && ({row_reg, col_reg}<18'b011000111010010111)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011000111010010111) && ({row_reg, col_reg}<18'b011000111010011100)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b011000111010011100)) color_data = 12'b010110101110;
		if(({row_reg, col_reg}==18'b011000111010011101)) color_data = 12'b011010111111;
		if(({row_reg, col_reg}>=18'b011000111010011110) && ({row_reg, col_reg}<18'b011000111010100000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011000111010100000)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b011000111010100001) && ({row_reg, col_reg}<18'b011000111010100101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011000111010100101) && ({row_reg, col_reg}<18'b011000111010101000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b011000111010101000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011000111010101001)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011000111010101010) && ({row_reg, col_reg}<18'b011000111010110010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011000111010110010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011000111010110011) && ({row_reg, col_reg}<18'b011000111011000001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011000111011000001)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011000111011000010) && ({row_reg, col_reg}<18'b011000111011001001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011000111011001001)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011000111011001010) && ({row_reg, col_reg}<18'b011000111011011010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011000111011011010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011000111011011011) && ({row_reg, col_reg}<18'b011000111011110011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011000111011110011)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011000111011110100) && ({row_reg, col_reg}<18'b011000111011110111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011000111011110111)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011000111011111000) && ({row_reg, col_reg}<18'b011000111011111110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011000111011111110) && ({row_reg, col_reg}<18'b011000111100000000)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b011000111100000000) && ({row_reg, col_reg}<18'b011001000000010010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011001000000010010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b011001000000010011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011001000000010100) && ({row_reg, col_reg}<18'b011001000000010110)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}==18'b011001000000010110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011001000000010111) && ({row_reg, col_reg}<18'b011001000000011001)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}>=18'b011001000000011001) && ({row_reg, col_reg}<18'b011001000000011011)) color_data = 12'b010110011111;
		if(({row_reg, col_reg}==18'b011001000000011011)) color_data = 12'b010010001110;
		if(({row_reg, col_reg}==18'b011001000000011100)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011001000000011101)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011001000000011110)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b011001000000011111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011001000000100000) && ({row_reg, col_reg}<18'b011001000000100011)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011001000000100011)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011001000000100100)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011001000000100101)) color_data = 12'b010010001110;
		if(({row_reg, col_reg}==18'b011001000000100110)) color_data = 12'b010010011110;
		if(({row_reg, col_reg}==18'b011001000000100111)) color_data = 12'b010010001110;
		if(({row_reg, col_reg}==18'b011001000000101000)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}==18'b011001000000101001)) color_data = 12'b010010001110;
		if(({row_reg, col_reg}>=18'b011001000000101010) && ({row_reg, col_reg}<18'b011001000000101100)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011001000000101100)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011001000000101101)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b011001000000101110)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011001000000101111) && ({row_reg, col_reg}<18'b011001000000110011)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011001000000110011) && ({row_reg, col_reg}<18'b011001000000110110)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011001000000110110)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011001000000110111)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011001000000111000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011001000000111001) && ({row_reg, col_reg}<18'b011001000000111100)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011001000000111100) && ({row_reg, col_reg}<18'b011001000000111111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011001000000111111)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011001000001000000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011001000001000001)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011001000001000010)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011001000001000011)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011001000001000100)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b011001000001000101)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011001000001000110)) color_data = 12'b010010011110;
		if(({row_reg, col_reg}==18'b011001000001000111)) color_data = 12'b010110101111;
		if(({row_reg, col_reg}==18'b011001000001001000)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==18'b011001000001001001)) color_data = 12'b010110101111;
		if(({row_reg, col_reg}==18'b011001000001001010)) color_data = 12'b010010011110;
		if(({row_reg, col_reg}==18'b011001000001001011)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==18'b011001000001001100)) color_data = 12'b010010011110;
		if(({row_reg, col_reg}>=18'b011001000001001101) && ({row_reg, col_reg}<18'b011001000001010000)) color_data = 12'b010110101110;
		if(({row_reg, col_reg}==18'b011001000001010000)) color_data = 12'b011011001111;
		if(({row_reg, col_reg}>=18'b011001000001010001) && ({row_reg, col_reg}<18'b011001000001011100)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}==18'b011001000001011100)) color_data = 12'b011111001111;
		if(({row_reg, col_reg}==18'b011001000001011101)) color_data = 12'b011011001111;
		if(({row_reg, col_reg}>=18'b011001000001011110) && ({row_reg, col_reg}<18'b011001000001100000)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b011001000001100000)) color_data = 12'b001010001101;
		if(({row_reg, col_reg}==18'b011001000001100001)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011001000001100010)) color_data = 12'b001110011101;
		if(({row_reg, col_reg}>=18'b011001000001100011) && ({row_reg, col_reg}<18'b011001000001100101)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}>=18'b011001000001100101) && ({row_reg, col_reg}<18'b011001000001100111)) color_data = 12'b011111011110;
		if(({row_reg, col_reg}==18'b011001000001100111)) color_data = 12'b100011101110;
		if(({row_reg, col_reg}>=18'b011001000001101000) && ({row_reg, col_reg}<18'b011001000001110110)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b011001000001110110)) color_data = 12'b011011011101;
		if(({row_reg, col_reg}==18'b011001000001110111)) color_data = 12'b011011011110;
		if(({row_reg, col_reg}>=18'b011001000001111000) && ({row_reg, col_reg}<18'b011001000001111010)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}==18'b011001000001111010)) color_data = 12'b011011001110;
		if(({row_reg, col_reg}==18'b011001000001111011)) color_data = 12'b010010101100;
		if(({row_reg, col_reg}==18'b011001000001111100)) color_data = 12'b001110011011;
		if(({row_reg, col_reg}==18'b011001000001111101)) color_data = 12'b010010101100;
		if(({row_reg, col_reg}==18'b011001000001111110)) color_data = 12'b010010101101;
		if(({row_reg, col_reg}==18'b011001000001111111)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b011001000010000000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011001000010000001)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b011001000010000010)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011001000010000011)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b011001000010000100)) color_data = 12'b011011001111;
		if(({row_reg, col_reg}>=18'b011001000010000101) && ({row_reg, col_reg}<18'b011001000010001001)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}>=18'b011001000010001001) && ({row_reg, col_reg}<18'b011001000010001011)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}>=18'b011001000010001011) && ({row_reg, col_reg}<18'b011001000010001101)) color_data = 12'b100011011111;
		if(({row_reg, col_reg}==18'b011001000010001101)) color_data = 12'b011111001111;
		if(({row_reg, col_reg}==18'b011001000010001110)) color_data = 12'b010010001100;
		if(({row_reg, col_reg}>=18'b011001000010001111) && ({row_reg, col_reg}<18'b011001000010010001)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}>=18'b011001000010010001) && ({row_reg, col_reg}<18'b011001000010010011)) color_data = 12'b010010001110;
		if(({row_reg, col_reg}>=18'b011001000010010011) && ({row_reg, col_reg}<18'b011001000010011100)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}==18'b011001000010011100)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011001000010011101)) color_data = 12'b011010111111;
		if(({row_reg, col_reg}>=18'b011001000010011110) && ({row_reg, col_reg}<18'b011001000010100011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011001000010100011)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b011001000010100100) && ({row_reg, col_reg}<18'b011001000010110000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011001000010110000) && ({row_reg, col_reg}<18'b011001000010110011)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011001000010110011) && ({row_reg, col_reg}<18'b011001000010111100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011001000010111100)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011001000010111101) && ({row_reg, col_reg}<18'b011001000011111101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011001000011111101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b011001000011111110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011001000011111111)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b011001000100000000) && ({row_reg, col_reg}<18'b011001001000001100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011001001000001100) && ({row_reg, col_reg}<18'b011001001000010000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011001001000010000) && ({row_reg, col_reg}<18'b011001001000010100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011001001000010100) && ({row_reg, col_reg}<18'b011001001000010110)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011001001000010110)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==18'b011001001000010111)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}>=18'b011001001000011000) && ({row_reg, col_reg}<18'b011001001000011011)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011001001000011011)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b011001001000011100) && ({row_reg, col_reg}<18'b011001001000011110)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011001001000011110)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b011001001000011111)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b011001001000100000)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011001001000100001)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b011001001000100010) && ({row_reg, col_reg}<18'b011001001000100100)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011001001000100100)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}==18'b011001001000100101)) color_data = 12'b010110011111;
		if(({row_reg, col_reg}==18'b011001001000100110)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b011001001000100111) && ({row_reg, col_reg}<18'b011001001000101001)) color_data = 12'b010110101111;
		if(({row_reg, col_reg}==18'b011001001000101001)) color_data = 12'b010110011111;
		if(({row_reg, col_reg}>=18'b011001001000101010) && ({row_reg, col_reg}<18'b011001001000101111)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011001001000101111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011001001000110000) && ({row_reg, col_reg}<18'b011001001000110010)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b011001001000110010)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}>=18'b011001001000110011) && ({row_reg, col_reg}<18'b011001001000111000)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b011001001000111000)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011001001000111001)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b011001001000111010)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011001001000111011) && ({row_reg, col_reg}<18'b011001001000111111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011001001000111111) && ({row_reg, col_reg}<18'b011001001001000010)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011001001001000010) && ({row_reg, col_reg}<18'b011001001001000100)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011001001001000100)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011001001001000101)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011001001001000110)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011001001001000111)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b011001001001001000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011001001001001001)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011001001001001010)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011001001001001011)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011001001001001100)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011001001001001101) && ({row_reg, col_reg}<18'b011001001001010001)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011001001001010001)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}>=18'b011001001001010010) && ({row_reg, col_reg}<18'b011001001001010100)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}>=18'b011001001001010100) && ({row_reg, col_reg}<18'b011001001001011100)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}>=18'b011001001001011100) && ({row_reg, col_reg}<18'b011001001001011110)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b011001001001011110)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b011001001001011111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011001001001100000)) color_data = 12'b001010001101;
		if(({row_reg, col_reg}==18'b011001001001100001)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011001001001100010)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011001001001100011)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b011001001001100100)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b011001001001100101)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b011001001001100110)) color_data = 12'b001110011010;
		if(({row_reg, col_reg}==18'b011001001001100111)) color_data = 12'b010110111100;
		if(({row_reg, col_reg}==18'b011001001001101000)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b011001001001101001)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b011001001001101010) && ({row_reg, col_reg}<18'b011001001001110100)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b011001001001110100)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b011001001001110101)) color_data = 12'b011111011110;
		if(({row_reg, col_reg}==18'b011001001001110110)) color_data = 12'b001110011010;
		if(({row_reg, col_reg}==18'b011001001001110111)) color_data = 12'b001010001010;
		if(({row_reg, col_reg}==18'b011001001001111000)) color_data = 12'b001110011011;
		if(({row_reg, col_reg}==18'b011001001001111001)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b011001001001111010)) color_data = 12'b010010101100;
		if(({row_reg, col_reg}==18'b011001001001111011)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b011001001001111100)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b011001001001111101)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b011001001001111110)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b011001001001111111)) color_data = 12'b010110111110;
		if(({row_reg, col_reg}==18'b011001001010000000)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}>=18'b011001001010000001) && ({row_reg, col_reg}<18'b011001001010000100)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011001001010000100)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b011001001010000101)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b011001001010000110)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b011001001010000111)) color_data = 12'b001010001011;
		if(({row_reg, col_reg}==18'b011001001010001000)) color_data = 12'b001110001011;
		if(({row_reg, col_reg}==18'b011001001010001001)) color_data = 12'b010110101101;
		if(({row_reg, col_reg}==18'b011001001010001010)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}>=18'b011001001010001011) && ({row_reg, col_reg}<18'b011001001010001101)) color_data = 12'b011010111101;
		if(({row_reg, col_reg}==18'b011001001010001101)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==18'b011001001010001110)) color_data = 12'b010110101110;
		if(({row_reg, col_reg}>=18'b011001001010001111) && ({row_reg, col_reg}<18'b011001001010011011)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011001001010011011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011001001010011100) && ({row_reg, col_reg}<18'b011001001010011110)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b011001001010011110) && ({row_reg, col_reg}<18'b011001001010111100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011001001010111100) && ({row_reg, col_reg}<18'b011001001010111110)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b011001001010111110) && ({row_reg, col_reg}<18'b011001010000001010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011001010000001010) && ({row_reg, col_reg}<18'b011001010000010000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011001010000010000) && ({row_reg, col_reg}<18'b011001010000010100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011001010000010100) && ({row_reg, col_reg}<18'b011001010000010110)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011001010000010110)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==18'b011001010000010111)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011001010000011000)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011001010000011001)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011001010000011010)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b011001010000011011)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011001010000011100) && ({row_reg, col_reg}<18'b011001010000011110)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011001010000011110)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b011001010000011111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011001010000100000) && ({row_reg, col_reg}<18'b011001010000100100)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011001010000100100)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}==18'b011001010000100101)) color_data = 12'b010110011111;
		if(({row_reg, col_reg}>=18'b011001010000100110) && ({row_reg, col_reg}<18'b011001010000101001)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011001010000101001)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}>=18'b011001010000101010) && ({row_reg, col_reg}<18'b011001010000110000)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011001010000110000) && ({row_reg, col_reg}<18'b011001010000110010)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b011001010000110010)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011001010000110011)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b011001010000110100)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b011001010000110101) && ({row_reg, col_reg}<18'b011001010000110111)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b011001010000110111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011001010000111000)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b011001010000111001) && ({row_reg, col_reg}<18'b011001010000111110)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b011001010000111110)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b011001010000111111)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011001010001000000) && ({row_reg, col_reg}<18'b011001010001000011)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011001010001000011) && ({row_reg, col_reg}<18'b011001010001001000)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011001010001001000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011001010001001001) && ({row_reg, col_reg}<18'b011001010001001011)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011001010001001011)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011001010001001100)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}==18'b011001010001001101)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011001010001001110)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011001010001001111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011001010001010000)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b011001010001010001) && ({row_reg, col_reg}<18'b011001010001010100)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011001010001010100)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b011001010001010101) && ({row_reg, col_reg}<18'b011001010001011001)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b011001010001011001)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011001010001011010)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b011001010001011011)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011001010001011100)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b011001010001011101)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011001010001011110)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011001010001011111)) color_data = 12'b001001101101;
		if(({row_reg, col_reg}==18'b011001010001100000)) color_data = 12'b001010001101;
		if(({row_reg, col_reg}==18'b011001010001100001)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}==18'b011001010001100010)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011001010001100011)) color_data = 12'b001010001101;
		if(({row_reg, col_reg}==18'b011001010001100100)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011001010001100101)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b011001010001100110)) color_data = 12'b000101111010;
		if(({row_reg, col_reg}==18'b011001010001100111)) color_data = 12'b010010101100;
		if(({row_reg, col_reg}>=18'b011001010001101000) && ({row_reg, col_reg}<18'b011001010001101010)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b011001010001101010) && ({row_reg, col_reg}<18'b011001010001110010)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b011001010001110010)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b011001010001110011) && ({row_reg, col_reg}<18'b011001010001110101)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b011001010001110101)) color_data = 12'b011111011110;
		if(({row_reg, col_reg}==18'b011001010001110110)) color_data = 12'b001010001010;
		if(({row_reg, col_reg}==18'b011001010001110111)) color_data = 12'b000101111010;
		if(({row_reg, col_reg}==18'b011001010001111000)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b011001010001111001)) color_data = 12'b000101111010;
		if(({row_reg, col_reg}==18'b011001010001111010)) color_data = 12'b010110111101;
		if(({row_reg, col_reg}==18'b011001010001111011)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b011001010001111100)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}>=18'b011001010001111101) && ({row_reg, col_reg}<18'b011001010001111111)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b011001010001111111)) color_data = 12'b010010111101;
		if(({row_reg, col_reg}>=18'b011001010010000000) && ({row_reg, col_reg}<18'b011001010010000010)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011001010010000010)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b011001010010000011)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011001010010000100) && ({row_reg, col_reg}<18'b011001010010000110)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011001010010000110)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b011001010010000111)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011001010010001000)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b011001010010001001)) color_data = 12'b010110101110;
		if(({row_reg, col_reg}==18'b011001010010001010)) color_data = 12'b011010111111;
		if(({row_reg, col_reg}==18'b011001010010001011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011001010010001100)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}==18'b011001010010001101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011001010010001110)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}==18'b011001010010001111)) color_data = 12'b011110111111;
		if(({row_reg, col_reg}>=18'b011001010010010000) && ({row_reg, col_reg}<18'b011001010010011101)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b011001010010011101) && ({row_reg, col_reg}<18'b011001010010101001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011001010010101001) && ({row_reg, col_reg}<18'b011001010010101100)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011001010010101100) && ({row_reg, col_reg}<18'b011001010010111100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011001010010111100) && ({row_reg, col_reg}<18'b011001010010111110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011001010010111110) && ({row_reg, col_reg}<18'b011001010011000000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011001010011000000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011001010011000001) && ({row_reg, col_reg}<18'b011001010011001010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011001010011001010)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b011001010011001011) && ({row_reg, col_reg}<18'b011001011000001011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011001011000001011) && ({row_reg, col_reg}<18'b011001011000010000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011001011000010000) && ({row_reg, col_reg}<18'b011001011000010100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011001011000010100) && ({row_reg, col_reg}<18'b011001011000010110)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011001011000010110)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}>=18'b011001011000010111) && ({row_reg, col_reg}<18'b011001011000011100)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011001011000011100)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}==18'b011001011000011101)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011001011000011110)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011001011000011111) && ({row_reg, col_reg}<18'b011001011000100100)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011001011000100100)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}==18'b011001011000100101)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}>=18'b011001011000100110) && ({row_reg, col_reg}<18'b011001011000101001)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011001011000101001)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}>=18'b011001011000101010) && ({row_reg, col_reg}<18'b011001011000101100)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}>=18'b011001011000101100) && ({row_reg, col_reg}<18'b011001011000110001)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011001011000110001)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b011001011000110010)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011001011000110011) && ({row_reg, col_reg}<18'b011001011000110110)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b011001011000110110)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b011001011000110111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011001011000111000) && ({row_reg, col_reg}<18'b011001011000111010)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b011001011000111010) && ({row_reg, col_reg}<18'b011001011000111110)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}>=18'b011001011000111110) && ({row_reg, col_reg}<18'b011001011001000000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011001011001000000) && ({row_reg, col_reg}<18'b011001011001000010)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b011001011001000010) && ({row_reg, col_reg}<18'b011001011001000111)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011001011001000111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011001011001001000)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011001011001001001) && ({row_reg, col_reg}<18'b011001011001001011)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b011001011001001011)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011001011001001100) && ({row_reg, col_reg}<18'b011001011001001111)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b011001011001001111)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}>=18'b011001011001010000) && ({row_reg, col_reg}<18'b011001011001010010)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b011001011001010010) && ({row_reg, col_reg}<18'b011001011001010110)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}>=18'b011001011001010110) && ({row_reg, col_reg}<18'b011001011001011000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011001011001011000)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}>=18'b011001011001011001) && ({row_reg, col_reg}<18'b011001011001011100)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011001011001011100)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011001011001011101)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011001011001011110)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b011001011001011111)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b011001011001100000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011001011001100001)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b011001011001100010)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011001011001100011)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}==18'b011001011001100100)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011001011001100101)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b011001011001100110)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b011001011001100111)) color_data = 12'b010110101101;
		if(({row_reg, col_reg}>=18'b011001011001101000) && ({row_reg, col_reg}<18'b011001011001101010)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b011001011001101010)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b011001011001101011) && ({row_reg, col_reg}<18'b011001011001101101)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b011001011001101101) && ({row_reg, col_reg}<18'b011001011001110000)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b011001011001110000) && ({row_reg, col_reg}<18'b011001011001110011)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b011001011001110011)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}==18'b011001011001110100)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b011001011001110101)) color_data = 12'b011111101111;
		if(({row_reg, col_reg}==18'b011001011001110110)) color_data = 12'b001010001010;
		if(({row_reg, col_reg}==18'b011001011001110111)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b011001011001111000)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b011001011001111001)) color_data = 12'b000101111011;
		if(({row_reg, col_reg}==18'b011001011001111010)) color_data = 12'b010110111110;
		if(({row_reg, col_reg}==18'b011001011001111011)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b011001011001111100)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}>=18'b011001011001111101) && ({row_reg, col_reg}<18'b011001011001111111)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b011001011001111111)) color_data = 12'b010110111101;
		if(({row_reg, col_reg}==18'b011001011010000000)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011001011010000001)) color_data = 12'b001010001101;
		if(({row_reg, col_reg}==18'b011001011010000010)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b011001011010000011)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011001011010000100)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011001011010000101)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011001011010000110)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011001011010000111)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011001011010001000)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}==18'b011001011010001001)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==18'b011001011010001010)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b011001011010001011) && ({row_reg, col_reg}<18'b011001011010010000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011001011010010000) && ({row_reg, col_reg}<18'b011001011010010011)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b011001011010010011) && ({row_reg, col_reg}<18'b011001011010011001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011001011010011001) && ({row_reg, col_reg}<18'b011001011010011100)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b011001011010011100) && ({row_reg, col_reg}<18'b011001011010100111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011001011010100111) && ({row_reg, col_reg}<18'b011001011010110101)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b011001011010110101) && ({row_reg, col_reg}<18'b011001100000001100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011001100000001100) && ({row_reg, col_reg}<18'b011001100000010000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011001100000010000) && ({row_reg, col_reg}<18'b011001100000010100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011001100000010100) && ({row_reg, col_reg}<18'b011001100000010110)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011001100000010110)) color_data = 12'b010010011110;
		if(({row_reg, col_reg}>=18'b011001100000010111) && ({row_reg, col_reg}<18'b011001100000011011)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011001100000011011)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011001100000011100) && ({row_reg, col_reg}<18'b011001100000011110)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011001100000011110)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011001100000011111) && ({row_reg, col_reg}<18'b011001100000100001)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011001100000100001) && ({row_reg, col_reg}<18'b011001100000100100)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b011001100000100100)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}==18'b011001100000100101)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==18'b011001100000100110)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011001100000100111)) color_data = 12'b011110111111;
		if(({row_reg, col_reg}==18'b011001100000101000)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011001100000101001)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}>=18'b011001100000101010) && ({row_reg, col_reg}<18'b011001100000110000)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}>=18'b011001100000110000) && ({row_reg, col_reg}<18'b011001100000110011)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011001100000110011)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011001100000110100)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011001100000110101) && ({row_reg, col_reg}<18'b011001100000111000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011001100000111000)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}>=18'b011001100000111001) && ({row_reg, col_reg}<18'b011001100000111011)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b011001100000111011) && ({row_reg, col_reg}<18'b011001100000111101)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}>=18'b011001100000111101) && ({row_reg, col_reg}<18'b011001100001000000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011001100001000000) && ({row_reg, col_reg}<18'b011001100001000010)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}>=18'b011001100001000010) && ({row_reg, col_reg}<18'b011001100001000101)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011001100001000101) && ({row_reg, col_reg}<18'b011001100001001000)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011001100001001000) && ({row_reg, col_reg}<18'b011001100001001010)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b011001100001001010) && ({row_reg, col_reg}<18'b011001100001001100)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011001100001001100) && ({row_reg, col_reg}<18'b011001100001001111)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b011001100001001111)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}>=18'b011001100001010000) && ({row_reg, col_reg}<18'b011001100001010010)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b011001100001010010) && ({row_reg, col_reg}<18'b011001100001011001)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}>=18'b011001100001011001) && ({row_reg, col_reg}<18'b011001100001011011)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b011001100001011011) && ({row_reg, col_reg}<18'b011001100001011101)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011001100001011101) && ({row_reg, col_reg}<18'b011001100001100001)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b011001100001100001)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}>=18'b011001100001100010) && ({row_reg, col_reg}<18'b011001100001100100)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b011001100001100100)) color_data = 12'b001001101101;
		if(({row_reg, col_reg}==18'b011001100001100101)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}==18'b011001100001100110)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b011001100001100111)) color_data = 12'b010110101110;
		if(({row_reg, col_reg}>=18'b011001100001101000) && ({row_reg, col_reg}<18'b011001100001101111)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b011001100001101111)) color_data = 12'b100011111111;
		if(({row_reg, col_reg}>=18'b011001100001110000) && ({row_reg, col_reg}<18'b011001100001110011)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}>=18'b011001100001110011) && ({row_reg, col_reg}<18'b011001100001110101)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b011001100001110101)) color_data = 12'b011111011111;
		if(({row_reg, col_reg}==18'b011001100001110110)) color_data = 12'b001110011100;
		if(({row_reg, col_reg}==18'b011001100001110111)) color_data = 12'b001010001100;
		if(({row_reg, col_reg}==18'b011001100001111000)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b011001100001111001)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011001100001111010)) color_data = 12'b010110101110;
		if(({row_reg, col_reg}==18'b011001100001111011)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b011001100001111100)) color_data = 12'b100111101111;
		if(({row_reg, col_reg}==18'b011001100001111101)) color_data = 12'b100111111111;
		if(({row_reg, col_reg}==18'b011001100001111110)) color_data = 12'b100011101111;
		if(({row_reg, col_reg}==18'b011001100001111111)) color_data = 12'b010110101110;
		if(({row_reg, col_reg}>=18'b011001100010000000) && ({row_reg, col_reg}<18'b011001100010000010)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b011001100010000010) && ({row_reg, col_reg}<18'b011001100010000100)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011001100010000100) && ({row_reg, col_reg}<18'b011001100010000110)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011001100010000110) && ({row_reg, col_reg}<18'b011001100010001000)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b011001100010001000)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}==18'b011001100010001001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011001100010001010)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b011001100010001011) && ({row_reg, col_reg}<18'b011001100010010111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011001100010010111)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011001100010011000) && ({row_reg, col_reg}<18'b011001100010100111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011001100010100111)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011001100010101000) && ({row_reg, col_reg}<18'b011001100010101010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011001100010101010) && ({row_reg, col_reg}<18'b011001100010110000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011001100010110000) && ({row_reg, col_reg}<18'b011001100010111001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011001100010111001)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b011001100010111010) && ({row_reg, col_reg}<18'b011001101000010001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011001101000010001)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011001101000010010) && ({row_reg, col_reg}<18'b011001101000010100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011001101000010100) && ({row_reg, col_reg}<18'b011001101000010110)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011001101000010110)) color_data = 12'b010010011110;
		if(({row_reg, col_reg}==18'b011001101000010111)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b011001101000011000)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011001101000011001) && ({row_reg, col_reg}<18'b011001101000011011)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011001101000011011)) color_data = 12'b010010001110;
		if(({row_reg, col_reg}>=18'b011001101000011100) && ({row_reg, col_reg}<18'b011001101000011110)) color_data = 12'b010110011111;
		if(({row_reg, col_reg}>=18'b011001101000011110) && ({row_reg, col_reg}<18'b011001101000100101)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}>=18'b011001101000100101) && ({row_reg, col_reg}<18'b011001101000101000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011001101000101000)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011001101000101001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011001101000101010)) color_data = 12'b010110011101;
		if(({row_reg, col_reg}>=18'b011001101000101011) && ({row_reg, col_reg}<18'b011001101000110000)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}>=18'b011001101000110000) && ({row_reg, col_reg}<18'b011001101000110011)) color_data = 12'b010110011111;
		if(({row_reg, col_reg}==18'b011001101000110011)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}==18'b011001101000110100)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b011001101000110101) && ({row_reg, col_reg}<18'b011001101000111001)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011001101000111001) && ({row_reg, col_reg}<18'b011001101000111011)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b011001101000111011)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b011001101000111100)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b011001101000111101)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b011001101000111110)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011001101000111111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011001101001000000) && ({row_reg, col_reg}<18'b011001101001000011)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b011001101001000011)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011001101001000100)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011001101001000101) && ({row_reg, col_reg}<18'b011001101001000111)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011001101001000111)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b011001101001001000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011001101001001001)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011001101001001010)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011001101001001011) && ({row_reg, col_reg}<18'b011001101001001111)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011001101001001111) && ({row_reg, col_reg}<18'b011001101001010010)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b011001101001010010) && ({row_reg, col_reg}<18'b011001101001011010)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b011001101001011010)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011001101001011011) && ({row_reg, col_reg}<18'b011001101001011101)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011001101001011101)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011001101001011110) && ({row_reg, col_reg}<18'b011001101001100100)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b011001101001100100)) color_data = 12'b001001101101;
		if(({row_reg, col_reg}==18'b011001101001100101)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011001101001100110)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011001101001100111)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b011001101001101000)) color_data = 12'b010110101110;
		if(({row_reg, col_reg}>=18'b011001101001101001) && ({row_reg, col_reg}<18'b011001101001101011)) color_data = 12'b010110101101;
		if(({row_reg, col_reg}>=18'b011001101001101011) && ({row_reg, col_reg}<18'b011001101001101101)) color_data = 12'b010010101101;
		if(({row_reg, col_reg}==18'b011001101001101101)) color_data = 12'b010110101101;
		if(({row_reg, col_reg}==18'b011001101001101110)) color_data = 12'b010110111101;
		if(({row_reg, col_reg}>=18'b011001101001101111) && ({row_reg, col_reg}<18'b011001101001110010)) color_data = 12'b010010101101;
		if(({row_reg, col_reg}==18'b011001101001110010)) color_data = 12'b010110101101;
		if(({row_reg, col_reg}==18'b011001101001110011)) color_data = 12'b010110111110;
		if(({row_reg, col_reg}>=18'b011001101001110100) && ({row_reg, col_reg}<18'b011001101001110110)) color_data = 12'b010110101110;
		if(({row_reg, col_reg}==18'b011001101001110110)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b011001101001110111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011001101001111000)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b011001101001111001)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011001101001111010)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b011001101001111011)) color_data = 12'b010110101110;
		if(({row_reg, col_reg}==18'b011001101001111100)) color_data = 12'b010010101101;
		if(({row_reg, col_reg}==18'b011001101001111101)) color_data = 12'b010110101110;
		if(({row_reg, col_reg}==18'b011001101001111110)) color_data = 12'b010110111111;
		if(({row_reg, col_reg}==18'b011001101001111111)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b011001101010000000)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011001101010000001)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}>=18'b011001101010000010) && ({row_reg, col_reg}<18'b011001101010000100)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011001101010000100)) color_data = 12'b010010011110;
		if(({row_reg, col_reg}>=18'b011001101010000101) && ({row_reg, col_reg}<18'b011001101010000111)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==18'b011001101010000111)) color_data = 12'b010110011101;
		if(({row_reg, col_reg}==18'b011001101010001000)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}>=18'b011001101010001001) && ({row_reg, col_reg}<18'b011001101010011001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011001101010011001) && ({row_reg, col_reg}<18'b011001101010011011)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011001101010011011) && ({row_reg, col_reg}<18'b011001101010011101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011001101010011101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011001101010011110) && ({row_reg, col_reg}<18'b011001101010101101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011001101010101101) && ({row_reg, col_reg}<18'b011001101010110000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011001101010110000) && ({row_reg, col_reg}<18'b011001101010110110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011001101010110110) && ({row_reg, col_reg}<18'b011001101010111000)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b011001101010111000) && ({row_reg, col_reg}<18'b011001110000010000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011001110000010000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011001110000010001) && ({row_reg, col_reg}<18'b011001110000010101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011001110000010101)) color_data = 12'b011010111111;
		if(({row_reg, col_reg}==18'b011001110000010110)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==18'b011001110000010111)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}>=18'b011001110000011000) && ({row_reg, col_reg}<18'b011001110000011011)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011001110000011011)) color_data = 12'b010110011111;
		if(({row_reg, col_reg}==18'b011001110000011100)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011001110000011101)) color_data = 12'b011010111111;
		if(({row_reg, col_reg}>=18'b011001110000011110) && ({row_reg, col_reg}<18'b011001110000100010)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011001110000100010)) color_data = 12'b011010111111;
		if(({row_reg, col_reg}>=18'b011001110000100011) && ({row_reg, col_reg}<18'b011001110000100110)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b011001110000100110) && ({row_reg, col_reg}<18'b011001110000101000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011001110000101000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b011001110000101001)) color_data = 12'b011110111111;
		if(({row_reg, col_reg}==18'b011001110000101010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011001110000101011)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}>=18'b011001110000101100) && ({row_reg, col_reg}<18'b011001110000110011)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011001110000110011)) color_data = 12'b010010001110;
		if(({row_reg, col_reg}==18'b011001110000110100)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b011001110000110101)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011001110000110110) && ({row_reg, col_reg}<18'b011001110000111000)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011001110000111000) && ({row_reg, col_reg}<18'b011001110000111011)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011001110000111011)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}>=18'b011001110000111100) && ({row_reg, col_reg}<18'b011001110000111110)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b011001110000111110) && ({row_reg, col_reg}<18'b011001110001000000)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011001110001000000) && ({row_reg, col_reg}<18'b011001110001000011)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011001110001000011)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011001110001000100) && ({row_reg, col_reg}<18'b011001110001000110)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011001110001000110) && ({row_reg, col_reg}<18'b011001110001001000)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b011001110001001000) && ({row_reg, col_reg}<18'b011001110001001110)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011001110001001110)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011001110001001111) && ({row_reg, col_reg}<18'b011001110001010001)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011001110001010001)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b011001110001010010)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011001110001010011)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011001110001010100) && ({row_reg, col_reg}<18'b011001110001011000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011001110001011000) && ({row_reg, col_reg}<18'b011001110001011011)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b011001110001011011) && ({row_reg, col_reg}<18'b011001110001011110)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011001110001011110) && ({row_reg, col_reg}<18'b011001110001100001)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b011001110001100001)) color_data = 12'b001101111111;
		if(({row_reg, col_reg}==18'b011001110001100010)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b011001110001100011)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}==18'b011001110001100100)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b011001110001100101)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}>=18'b011001110001100110) && ({row_reg, col_reg}<18'b011001110001101001)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011001110001101001)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}>=18'b011001110001101010) && ({row_reg, col_reg}<18'b011001110001101101)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b011001110001101101) && ({row_reg, col_reg}<18'b011001110001110001)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}>=18'b011001110001110001) && ({row_reg, col_reg}<18'b011001110001110100)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011001110001110100)) color_data = 12'b000101101011;
		if(({row_reg, col_reg}>=18'b011001110001110101) && ({row_reg, col_reg}<18'b011001110001110111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011001110001110111)) color_data = 12'b000101101101;
		if(({row_reg, col_reg}==18'b011001110001111000)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b011001110001111001)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011001110001111010)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}==18'b011001110001111011)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011001110001111100)) color_data = 12'b001001111011;
		if(({row_reg, col_reg}==18'b011001110001111101)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b011001110001111110) && ({row_reg, col_reg}<18'b011001110010000000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011001110010000000)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b011001110010000001)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b011001110010000010)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011001110010000011)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011001110010000100)) color_data = 12'b010110011111;
		if(({row_reg, col_reg}>=18'b011001110010000101) && ({row_reg, col_reg}<18'b011001110010000111)) color_data = 12'b011110111111;
		if(({row_reg, col_reg}==18'b011001110010000111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011001110010001000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b011001110010001001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011001110010001010)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}>=18'b011001110010001011) && ({row_reg, col_reg}<18'b011001110010010111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011001110010010111)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011001110010011000) && ({row_reg, col_reg}<18'b011001110010101101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011001110010101101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b011001110010101110)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}>=18'b011001110010101111) && ({row_reg, col_reg}<18'b011001110010110101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011001110010110101) && ({row_reg, col_reg}<18'b011001110010111001)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b011001110010111001) && ({row_reg, col_reg}<18'b011001111000010000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011001111000010000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011001111000010001) && ({row_reg, col_reg}<18'b011001111000010101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011001111000010101)) color_data = 12'b011010111111;
		if(({row_reg, col_reg}==18'b011001111000010110)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}>=18'b011001111000010111) && ({row_reg, col_reg}<18'b011001111000011011)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011001111000011011)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}>=18'b011001111000011100) && ({row_reg, col_reg}<18'b011001111000100100)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011001111000100100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011001111000100101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b011001111000100110)) color_data = 12'b011110111110;
		if(({row_reg, col_reg}>=18'b011001111000100111) && ({row_reg, col_reg}<18'b011001111000101010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011001111000101010) && ({row_reg, col_reg}<18'b011001111000101101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011001111000101101) && ({row_reg, col_reg}<18'b011001111000110000)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011001111000110000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011001111000110001) && ({row_reg, col_reg}<18'b011001111000110011)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011001111000110011)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}==18'b011001111000110100)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011001111000110101)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011001111000110110) && ({row_reg, col_reg}<18'b011001111000111000)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b011001111000111000)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011001111000111001) && ({row_reg, col_reg}<18'b011001111000111101)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011001111000111101) && ({row_reg, col_reg}<18'b011001111001000010)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011001111001000010)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011001111001000011)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011001111001000100) && ({row_reg, col_reg}<18'b011001111001000111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011001111001000111)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b011001111001001000)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b011001111001001001)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011001111001001010) && ({row_reg, col_reg}<18'b011001111001001101)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b011001111001001101)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011001111001001110)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011001111001001111)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011001111001010000) && ({row_reg, col_reg}<18'b011001111001010011)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011001111001010011) && ({row_reg, col_reg}<18'b011001111001010101)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}>=18'b011001111001010101) && ({row_reg, col_reg}<18'b011001111001010111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011001111001010111)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011001111001011000) && ({row_reg, col_reg}<18'b011001111001011010)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b011001111001011010) && ({row_reg, col_reg}<18'b011001111001011110)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011001111001011110) && ({row_reg, col_reg}<18'b011001111001100000)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b011001111001100000)) color_data = 12'b001101111111;
		if(({row_reg, col_reg}>=18'b011001111001100001) && ({row_reg, col_reg}<18'b011001111001100011)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b011001111001100011)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b011001111001100100)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011001111001100101)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b011001111001100110)) color_data = 12'b001010001101;
		if(({row_reg, col_reg}>=18'b011001111001100111) && ({row_reg, col_reg}<18'b011001111001101010)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011001111001101010)) color_data = 12'b001010001101;
		if(({row_reg, col_reg}>=18'b011001111001101011) && ({row_reg, col_reg}<18'b011001111001101101)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}>=18'b011001111001101101) && ({row_reg, col_reg}<18'b011001111001101111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011001111001101111)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011001111001110000)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b011001111001110001)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011001111001110010)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011001111001110011)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b011001111001110100)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b011001111001110101) && ({row_reg, col_reg}<18'b011001111001110111)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}==18'b011001111001110111)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b011001111001111000)) color_data = 12'b001101111111;
		if(({row_reg, col_reg}==18'b011001111001111001)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b011001111001111010)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}==18'b011001111001111011)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011001111001111100) && ({row_reg, col_reg}<18'b011001111001111110)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}>=18'b011001111001111110) && ({row_reg, col_reg}<18'b011001111010000000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011001111010000000)) color_data = 12'b001101111111;
		if(({row_reg, col_reg}==18'b011001111010000001)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b011001111010000010)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011001111010000011)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011001111010000100)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==18'b011001111010000101)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011001111010000110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011001111010000111)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}==18'b011001111010001000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011001111010001001)) color_data = 12'b011110111110;
		if(({row_reg, col_reg}>=18'b011001111010001010) && ({row_reg, col_reg}<18'b011001111010001101)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}>=18'b011001111010001101) && ({row_reg, col_reg}<18'b011001111010001111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011001111010001111) && ({row_reg, col_reg}<18'b011001111010010001)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b011001111010010001) && ({row_reg, col_reg}<18'b011001111010010101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011001111010010101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011001111010010110) && ({row_reg, col_reg}<18'b011001111010011000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011001111010011000) && ({row_reg, col_reg}<18'b011001111010100000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011001111010100000) && ({row_reg, col_reg}<18'b011001111010110101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011001111010110101) && ({row_reg, col_reg}<18'b011001111010111010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011001111010111010) && ({row_reg, col_reg}<18'b011001111011000000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011001111011000000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011001111011000001) && ({row_reg, col_reg}<18'b011001111011000100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011001111011000100) && ({row_reg, col_reg}<18'b011001111011000110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011001111011000110) && ({row_reg, col_reg}<18'b011001111011111011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011001111011111011)) color_data = 12'b011010101111;

		if(({row_reg, col_reg}>=18'b011001111011111100) && ({row_reg, col_reg}<18'b011010000000010000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011010000000010000) && ({row_reg, col_reg}<18'b011010000000010010)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}>=18'b011010000000010010) && ({row_reg, col_reg}<18'b011010000000010101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011010000000010101)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011010000000010110)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}>=18'b011010000000010111) && ({row_reg, col_reg}<18'b011010000000011010)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b011010000000011010)) color_data = 12'b001001101011;
		if(({row_reg, col_reg}==18'b011010000000011011)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==18'b011010000000011100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011010000000011101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b011010000000011110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011010000000011111)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011010000000100000) && ({row_reg, col_reg}<18'b011010000000100011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011010000000100011)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011010000000100100) && ({row_reg, col_reg}<18'b011010000000100110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011010000000100110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011010000000100111) && ({row_reg, col_reg}<18'b011010000000101001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011010000000101001)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b011010000000101010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011010000000101011) && ({row_reg, col_reg}<18'b011010000000101101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b011010000000101101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011010000000101110) && ({row_reg, col_reg}<18'b011010000000110000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011010000000110000) && ({row_reg, col_reg}<18'b011010000000110010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011010000000110010)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011010000000110011)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}>=18'b011010000000110100) && ({row_reg, col_reg}<18'b011010000000110111)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b011010000000110111)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011010000000111000)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011010000000111001)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011010000000111010)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b011010000000111011) && ({row_reg, col_reg}<18'b011010000000111111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011010000000111111)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011010000001000000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011010000001000001)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b011010000001000010)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011010000001000011)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}>=18'b011010000001000100) && ({row_reg, col_reg}<18'b011010000001001000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011010000001001000) && ({row_reg, col_reg}<18'b011010000001001101)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b011010000001001101) && ({row_reg, col_reg}<18'b011010000001010001)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011010000001010001)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011010000001010010)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b011010000001010011)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011010000001010100) && ({row_reg, col_reg}<18'b011010000001011000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011010000001011000) && ({row_reg, col_reg}<18'b011010000001011100)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b011010000001011100) && ({row_reg, col_reg}<18'b011010000001100000)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b011010000001100000)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011010000001100001)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b011010000001100010)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b011010000001100011) && ({row_reg, col_reg}<18'b011010000001100101)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011010000001100101) && ({row_reg, col_reg}<18'b011010000001101000)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}>=18'b011010000001101000) && ({row_reg, col_reg}<18'b011010000001101010)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011010000001101010)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011010000001101011)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011010000001101100) && ({row_reg, col_reg}<18'b011010000001101110)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011010000001101110) && ({row_reg, col_reg}<18'b011010000001110000)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b011010000001110000) && ({row_reg, col_reg}<18'b011010000001110010)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b011010000001110010)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011010000001110011)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b011010000001110100)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011010000001110101) && ({row_reg, col_reg}<18'b011010000001110111)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011010000001110111) && ({row_reg, col_reg}<18'b011010000001111100)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b011010000001111100) && ({row_reg, col_reg}<18'b011010000010000000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011010000010000000) && ({row_reg, col_reg}<18'b011010000010000010)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011010000010000010) && ({row_reg, col_reg}<18'b011010000010000100)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b011010000010000100)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}>=18'b011010000010000101) && ({row_reg, col_reg}<18'b011010000010001000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011010000010001000) && ({row_reg, col_reg}<18'b011010000010001010)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b011010000010001010) && ({row_reg, col_reg}<18'b011010001000010000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011010001000010000)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}==18'b011010001000010001)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011010001000010010) && ({row_reg, col_reg}<18'b011010001000010101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011010001000010101)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011010001000010110)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}>=18'b011010001000010111) && ({row_reg, col_reg}<18'b011010001000011010)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}==18'b011010001000011010)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b011010001000011011)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}>=18'b011010001000011100) && ({row_reg, col_reg}<18'b011010001000011110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011010001000011110)) color_data = 12'b011010101101;
		if(({row_reg, col_reg}>=18'b011010001000011111) && ({row_reg, col_reg}<18'b011010001000100010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011010001000100010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b011010001000100011)) color_data = 12'b011110111110;
		if(({row_reg, col_reg}==18'b011010001000100100)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011010001000100101) && ({row_reg, col_reg}<18'b011010001000101001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011010001000101001)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011010001000101010) && ({row_reg, col_reg}<18'b011010001000101100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011010001000101100)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011010001000101101) && ({row_reg, col_reg}<18'b011010001000110010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011010001000110010)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011010001000110011)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}==18'b011010001000110100)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011010001000110101)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b011010001000110110)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011010001000110111)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011010001000111000) && ({row_reg, col_reg}<18'b011010001000111011)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b011010001000111011)) color_data = 12'b010010011110;
		if(({row_reg, col_reg}==18'b011010001000111100)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}==18'b011010001000111101)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011010001000111110) && ({row_reg, col_reg}<18'b011010001001000000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011010001001000000) && ({row_reg, col_reg}<18'b011010001001000010)) color_data = 12'b001001111110;
		if(({row_reg, col_reg}==18'b011010001001000010)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011010001001000011)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}>=18'b011010001001000100) && ({row_reg, col_reg}<18'b011010001001000110)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011010001001000110) && ({row_reg, col_reg}<18'b011010001001001110)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b011010001001001110)) color_data = 12'b010010001110;
		if(({row_reg, col_reg}==18'b011010001001001111)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b011010001001010000) && ({row_reg, col_reg}<18'b011010001001010011)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011010001001010011)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011010001001010100)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011010001001010101)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}==18'b011010001001010110)) color_data = 12'b010010001110;
		if(({row_reg, col_reg}>=18'b011010001001010111) && ({row_reg, col_reg}<18'b011010001001011011)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}>=18'b011010001001011011) && ({row_reg, col_reg}<18'b011010001001100001)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}>=18'b011010001001100001) && ({row_reg, col_reg}<18'b011010001001100011)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b011010001001100011)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011010001001100100)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}==18'b011010001001100101)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b011010001001100110)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}==18'b011010001001100111)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b011010001001101000) && ({row_reg, col_reg}<18'b011010001001101101)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011010001001101101) && ({row_reg, col_reg}<18'b011010001001110000)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011010001001110000)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}>=18'b011010001001110001) && ({row_reg, col_reg}<18'b011010001001110011)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}>=18'b011010001001110011) && ({row_reg, col_reg}<18'b011010001001111100)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b011010001001111100)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}>=18'b011010001001111101) && ({row_reg, col_reg}<18'b011010001010000000)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}>=18'b011010001010000000) && ({row_reg, col_reg}<18'b011010001010000010)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011010001010000010)) color_data = 12'b010001111101;
		if(({row_reg, col_reg}==18'b011010001010000011)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}==18'b011010001010000100)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==18'b011010001010000101)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011010001010000110)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}>=18'b011010001010000111) && ({row_reg, col_reg}<18'b011010001010001001)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b011010001010001001) && ({row_reg, col_reg}<18'b011010010000010101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011010010000010101)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011010010000010110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011010010000010111)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}>=18'b011010010000011000) && ({row_reg, col_reg}<18'b011010010000011010)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b011010010000011010) && ({row_reg, col_reg}<18'b011010010000011101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011010010000011101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b011010010000011110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011010010000011111) && ({row_reg, col_reg}<18'b011010010000100001)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011010010000100001) && ({row_reg, col_reg}<18'b011010010000100110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011010010000100110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011010010000100111) && ({row_reg, col_reg}<18'b011010010000101001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011010010000101001)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011010010000101010) && ({row_reg, col_reg}<18'b011010010000101100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011010010000101100)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011010010000101101) && ({row_reg, col_reg}<18'b011010010000110010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011010010000110010)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011010010000110011)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b011010010000110100)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}>=18'b011010010000110101) && ({row_reg, col_reg}<18'b011010010000110111)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b011010010000110111)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b011010010000111000)) color_data = 12'b010110011111;
		if(({row_reg, col_reg}>=18'b011010010000111001) && ({row_reg, col_reg}<18'b011010010000111100)) color_data = 12'b010110101111;
		if(({row_reg, col_reg}==18'b011010010000111100)) color_data = 12'b010010011110;
		if(({row_reg, col_reg}==18'b011010010000111101)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}==18'b011010010000111110)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011010010000111111) && ({row_reg, col_reg}<18'b011010010001000011)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011010010001000011)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b011010010001000100)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011010010001000101)) color_data = 12'b001110001110;
		if(({row_reg, col_reg}==18'b011010010001000110)) color_data = 12'b010010011111;
		if(({row_reg, col_reg}==18'b011010010001000111)) color_data = 12'b010110101111;
		if(({row_reg, col_reg}>=18'b011010010001001000) && ({row_reg, col_reg}<18'b011010010001001111)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011010010001001111)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}>=18'b011010010001010000) && ({row_reg, col_reg}<18'b011010010001010100)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011010010001010100)) color_data = 12'b010010001110;
		if(({row_reg, col_reg}==18'b011010010001010101)) color_data = 12'b010110101111;
		if(({row_reg, col_reg}>=18'b011010010001010110) && ({row_reg, col_reg}<18'b011010010001011000)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011010010001011000)) color_data = 12'b010110101111;
		if(({row_reg, col_reg}>=18'b011010010001011001) && ({row_reg, col_reg}<18'b011010010001100010)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011010010001100010)) color_data = 12'b010110101111;
		if(({row_reg, col_reg}==18'b011010010001100011)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011010010001100100) && ({row_reg, col_reg}<18'b011010010001100110)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011010010001100110)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011010010001100111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011010010001101000)) color_data = 12'b001101111110;
		if(({row_reg, col_reg}==18'b011010010001101001)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011010010001101010) && ({row_reg, col_reg}<18'b011010010001101100)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011010010001101100) && ({row_reg, col_reg}<18'b011010010001101110)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011010010001101110) && ({row_reg, col_reg}<18'b011010010001110000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011010010001110000)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b011010010001110001)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==18'b011010010001110010)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011010010001110011)) color_data = 12'b010110101111;
		if(({row_reg, col_reg}>=18'b011010010001110100) && ({row_reg, col_reg}<18'b011010010001110110)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011010010001110110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011010010001110111) && ({row_reg, col_reg}<18'b011010010001111010)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011010010001111010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011010010001111011) && ({row_reg, col_reg}<18'b011010010010000100)) color_data = 12'b011010101111;

		if(({row_reg, col_reg}>=18'b011010010010000100) && ({row_reg, col_reg}<18'b011010011000010101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011010011000010101) && ({row_reg, col_reg}<18'b011010011000010111)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011010011000010111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011010011000011000) && ({row_reg, col_reg}<18'b011010011000011011)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b011010011000011011) && ({row_reg, col_reg}<18'b011010011000100011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011010011000100011)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011010011000100100) && ({row_reg, col_reg}<18'b011010011000100110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011010011000100110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011010011000100111) && ({row_reg, col_reg}<18'b011010011000110001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011010011000110001) && ({row_reg, col_reg}<18'b011010011000110011)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011010011000110011)) color_data = 12'b001110001100;
		if(({row_reg, col_reg}==18'b011010011000110100)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b011010011000110101)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b011010011000110110)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011010011000110111)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b011010011000111000)) color_data = 12'b010110101111;
		if(({row_reg, col_reg}>=18'b011010011000111001) && ({row_reg, col_reg}<18'b011010011000111100)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011010011000111100)) color_data = 12'b010010011110;
		if(({row_reg, col_reg}>=18'b011010011000111101) && ({row_reg, col_reg}<18'b011010011001000101)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011010011001000101)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b011010011001000110)) color_data = 12'b010110011111;
		if(({row_reg, col_reg}==18'b011010011001000111)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011010011001001000)) color_data = 12'b011010111111;
		if(({row_reg, col_reg}>=18'b011010011001001001) && ({row_reg, col_reg}<18'b011010011001001101)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011010011001001101)) color_data = 12'b011010111111;
		if(({row_reg, col_reg}==18'b011010011001001110)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011010011001001111)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==18'b011010011001010000)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b011010011001010001)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011010011001010010) && ({row_reg, col_reg}<18'b011010011001010100)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b011010011001010100)) color_data = 12'b010010011110;
		if(({row_reg, col_reg}>=18'b011010011001010101) && ({row_reg, col_reg}<18'b011010011001011011)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b011010011001011011) && ({row_reg, col_reg}<18'b011010011001011110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011010011001011110) && ({row_reg, col_reg}<18'b011010011001100000)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011010011001100000)) color_data = 12'b011010111111;
		if(({row_reg, col_reg}>=18'b011010011001100001) && ({row_reg, col_reg}<18'b011010011001100011)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011010011001100011)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}>=18'b011010011001100100) && ({row_reg, col_reg}<18'b011010011001101000)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011010011001101000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011010011001101001)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011010011001101010) && ({row_reg, col_reg}<18'b011010011001101100)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011010011001101100) && ({row_reg, col_reg}<18'b011010011001101110)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011010011001101110) && ({row_reg, col_reg}<18'b011010011001110000)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011010011001110000)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}==18'b011010011001110001)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==18'b011010011001110010)) color_data = 12'b011010111111;
		if(({row_reg, col_reg}>=18'b011010011001110011) && ({row_reg, col_reg}<18'b011010011001110101)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b011010011001110101) && ({row_reg, col_reg}<18'b011010011001111111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011010011001111111) && ({row_reg, col_reg}<18'b011010011010000100)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b011010011010000100) && ({row_reg, col_reg}<18'b011010011010000110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011010011010000110)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b011010011010000111) && ({row_reg, col_reg}<18'b011010100000010000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011010100000010000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011010100000010001) && ({row_reg, col_reg}<18'b011010100000100000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011010100000100000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011010100000100001) && ({row_reg, col_reg}<18'b011010100000100011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011010100000100011)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011010100000100100) && ({row_reg, col_reg}<18'b011010100000110001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011010100000110001) && ({row_reg, col_reg}<18'b011010100000110011)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011010100000110011)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}>=18'b011010100000110100) && ({row_reg, col_reg}<18'b011010100000110111)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b011010100000110111)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}==18'b011010100000111000)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b011010100000111001) && ({row_reg, col_reg}<18'b011010100000111100)) color_data = 12'b011010111111;
		if(({row_reg, col_reg}==18'b011010100000111100)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}>=18'b011010100000111101) && ({row_reg, col_reg}<18'b011010100001000010)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011010100001000010)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011010100001000011)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011010100001000100)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}==18'b011010100001000101)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011010100001000110)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}>=18'b011010100001000111) && ({row_reg, col_reg}<18'b011010100001001001)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b011010100001001001) && ({row_reg, col_reg}<18'b011010100001001101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011010100001001101) && ({row_reg, col_reg}<18'b011010100001001111)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011010100001001111)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==18'b011010100001010000)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b011010100001010001)) color_data = 12'b001001111100;
		if(({row_reg, col_reg}>=18'b011010100001010010) && ({row_reg, col_reg}<18'b011010100001010100)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b011010100001010100)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}>=18'b011010100001010101) && ({row_reg, col_reg}<18'b011010100001010111)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b011010100001010111) && ({row_reg, col_reg}<18'b011010100001011011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011010100001011011)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011010100001011100) && ({row_reg, col_reg}<18'b011010100001011111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011010100001011111)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011010100001100000) && ({row_reg, col_reg}<18'b011010100001100011)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011010100001100011)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}>=18'b011010100001100100) && ({row_reg, col_reg}<18'b011010100001101010)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011010100001101010) && ({row_reg, col_reg}<18'b011010100001101100)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}>=18'b011010100001101100) && ({row_reg, col_reg}<18'b011010100001110000)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011010100001110000)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}==18'b011010100001110001)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==18'b011010100001110010)) color_data = 12'b011110111111;
		if(({row_reg, col_reg}==18'b011010100001110011)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b011010100001110100) && ({row_reg, col_reg}<18'b011010100001110110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011010100001110110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011010100001110111) && ({row_reg, col_reg}<18'b011010100010000000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011010100010000000)) color_data = 12'b011010101111;

		if(({row_reg, col_reg}>=18'b011010100010000001) && ({row_reg, col_reg}<18'b011010101000100001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011010101000100001) && ({row_reg, col_reg}<18'b011010101000100011)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011010101000100011) && ({row_reg, col_reg}<18'b011010101000100110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011010101000100110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011010101000100111) && ({row_reg, col_reg}<18'b011010101000110000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011010101000110000) && ({row_reg, col_reg}<18'b011010101000110011)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011010101000110011)) color_data = 12'b010010001100;
		if(({row_reg, col_reg}>=18'b011010101000110100) && ({row_reg, col_reg}<18'b011010101000110111)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b011010101000110111)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}==18'b011010101000111000)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}>=18'b011010101000111001) && ({row_reg, col_reg}<18'b011010101000111100)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011010101000111100)) color_data = 12'b010010011101;
		if(({row_reg, col_reg}==18'b011010101000111101)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}>=18'b011010101000111110) && ({row_reg, col_reg}<18'b011010101001000010)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}>=18'b011010101001000010) && ({row_reg, col_reg}<18'b011010101001000101)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011010101001000101)) color_data = 12'b010010001101;
		if(({row_reg, col_reg}==18'b011010101001000110)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}>=18'b011010101001000111) && ({row_reg, col_reg}<18'b011010101001001001)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b011010101001001001) && ({row_reg, col_reg}<18'b011010101001001111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011010101001001111)) color_data = 12'b010110011101;
		if(({row_reg, col_reg}==18'b011010101001010000)) color_data = 12'b001110001101;
		if(({row_reg, col_reg}>=18'b011010101001010001) && ({row_reg, col_reg}<18'b011010101001010100)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}==18'b011010101001010100)) color_data = 12'b010010011101;
		if(({row_reg, col_reg}==18'b011010101001010101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011010101001010110)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011010101001010111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011010101001011000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011010101001011001) && ({row_reg, col_reg}<18'b011010101001011011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011010101001011011)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011010101001011100) && ({row_reg, col_reg}<18'b011010101001011111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011010101001011111)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b011010101001100000)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b011010101001100001) && ({row_reg, col_reg}<18'b011010101001100011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011010101001100011) && ({row_reg, col_reg}<18'b011010101001100110)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}>=18'b011010101001100110) && ({row_reg, col_reg}<18'b011010101001101011)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011010101001101011)) color_data = 12'b001101111100;
		if(({row_reg, col_reg}>=18'b011010101001101100) && ({row_reg, col_reg}<18'b011010101001101111)) color_data = 12'b001101111101;
		if(({row_reg, col_reg}==18'b011010101001101111)) color_data = 12'b001001111101;
		if(({row_reg, col_reg}==18'b011010101001110000)) color_data = 12'b010001111100;
		if(({row_reg, col_reg}==18'b011010101001110001)) color_data = 12'b010110011101;
		if(({row_reg, col_reg}>=18'b011010101001110010) && ({row_reg, col_reg}<18'b011010101001110110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011010101001110110)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b011010101001110111) && ({row_reg, col_reg}<18'b011010110000011110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011010110000011110) && ({row_reg, col_reg}<18'b011010110000100001)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011010110000100001) && ({row_reg, col_reg}<18'b011010110000100100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011010110000100100)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011010110000100101) && ({row_reg, col_reg}<18'b011010110000100111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011010110000100111)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011010110000101000) && ({row_reg, col_reg}<18'b011010110000110000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011010110000110000) && ({row_reg, col_reg}<18'b011010110000110011)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b011010110000110011) && ({row_reg, col_reg}<18'b011010110000110101)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}>=18'b011010110000110101) && ({row_reg, col_reg}<18'b011010110000110111)) color_data = 12'b010110011101;
		if(({row_reg, col_reg}==18'b011010110000110111)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}>=18'b011010110000111000) && ({row_reg, col_reg}<18'b011010110000111011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011010110000111011)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011010110000111100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011010110000111101) && ({row_reg, col_reg}<18'b011010110001000100)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==18'b011010110001000100)) color_data = 12'b010010011110;
		if(({row_reg, col_reg}==18'b011010110001000101)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==18'b011010110001000110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011010110001000111)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b011010110001001000) && ({row_reg, col_reg}<18'b011010110001001101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011010110001001101) && ({row_reg, col_reg}<18'b011010110001001111)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b011010110001001111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011010110001010000)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==18'b011010110001010001)) color_data = 12'b010110011101;
		if(({row_reg, col_reg}==18'b011010110001010010)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==18'b011010110001010011)) color_data = 12'b010110011101;
		if(({row_reg, col_reg}==18'b011010110001010100)) color_data = 12'b010110101110;
		if(({row_reg, col_reg}>=18'b011010110001010101) && ({row_reg, col_reg}<18'b011010110001010111)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011010110001010111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011010110001011000) && ({row_reg, col_reg}<18'b011010110001011110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b011010110001011110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011010110001011111)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b011010110001100000)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}>=18'b011010110001100001) && ({row_reg, col_reg}<18'b011010110001100011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011010110001100011)) color_data = 12'b010110011101;
		if(({row_reg, col_reg}>=18'b011010110001100100) && ({row_reg, col_reg}<18'b011010110001101111)) color_data = 12'b010110011110;
		if(({row_reg, col_reg}==18'b011010110001101111)) color_data = 12'b010010011110;
		if(({row_reg, col_reg}==18'b011010110001110000)) color_data = 12'b010110011101;

		if(({row_reg, col_reg}>=18'b011010110001110001) && ({row_reg, col_reg}<18'b011010111000011001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011010111000011001)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b011010111000011010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011010111000011011)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011010111000011100) && ({row_reg, col_reg}<18'b011010111000110000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011010111000110000) && ({row_reg, col_reg}<18'b011010111000110100)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011010111000110100)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}>=18'b011010111000110101) && ({row_reg, col_reg}<18'b011010111000111000)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b011010111000111000) && ({row_reg, col_reg}<18'b011010111000111010)) color_data = 12'b011110111111;
		if(({row_reg, col_reg}==18'b011010111000111010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011010111000111011)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}==18'b011010111000111100)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b011010111000111101) && ({row_reg, col_reg}<18'b011010111001000000)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}>=18'b011010111001000000) && ({row_reg, col_reg}<18'b011010111001000010)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011010111001000010)) color_data = 12'b011110111111;
		if(({row_reg, col_reg}>=18'b011010111001000011) && ({row_reg, col_reg}<18'b011010111001000111)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011010111001000111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011010111001001000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b011010111001001001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011010111001001010) && ({row_reg, col_reg}<18'b011010111001001111)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011010111001001111) && ({row_reg, col_reg}<18'b011010111001010001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011010111001010001) && ({row_reg, col_reg}<18'b011010111001010011)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011010111001010011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011010111001010100) && ({row_reg, col_reg}<18'b011010111001010110)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011010111001010110)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}>=18'b011010111001010111) && ({row_reg, col_reg}<18'b011010111001011001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011010111001011001) && ({row_reg, col_reg}<18'b011010111001011101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011010111001011101) && ({row_reg, col_reg}<18'b011010111001011111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011010111001011111)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b011010111001100000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011010111001100001)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}==18'b011010111001100010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011010111001100011)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}==18'b011010111001100100)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b011010111001100101) && ({row_reg, col_reg}<18'b011010111001100111)) color_data = 12'b011110101111;
		if(({row_reg, col_reg}>=18'b011010111001100111) && ({row_reg, col_reg}<18'b011010111001101001)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011010111001101001)) color_data = 12'b011010111111;
		if(({row_reg, col_reg}>=18'b011010111001101010) && ({row_reg, col_reg}<18'b011010111001110010)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011010111001110010)) color_data = 12'b011110111111;
		if(({row_reg, col_reg}>=18'b011010111001110011) && ({row_reg, col_reg}<18'b011010111010000010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011010111010000010)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b011010111010000011) && ({row_reg, col_reg}<18'b011011000000110101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011011000000110101)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b011011000000110110) && ({row_reg, col_reg}<18'b011011000000111111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011011000000111111) && ({row_reg, col_reg}<18'b011011000001000110)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b011011000001000110) && ({row_reg, col_reg}<18'b011011000001001010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011011000001001010) && ({row_reg, col_reg}<18'b011011000001001101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011011000001001101) && ({row_reg, col_reg}<18'b011011000001010001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011011000001010001)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}==18'b011011000001010010)) color_data = 12'b011010111111;
		if(({row_reg, col_reg}==18'b011011000001010011)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b011011000001010100) && ({row_reg, col_reg}<18'b011011000001011001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011011000001011001) && ({row_reg, col_reg}<18'b011011000001011101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011011000001011101) && ({row_reg, col_reg}<18'b011011000001100100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011011000001100100) && ({row_reg, col_reg}<18'b011011000001110000)) color_data = 12'b011010101111;

		if(({row_reg, col_reg}>=18'b011011000001110000) && ({row_reg, col_reg}<18'b011011001000110010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011011001000110010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011011001000110011) && ({row_reg, col_reg}<18'b011011001000110101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011011001000110101) && ({row_reg, col_reg}<18'b011011001000111000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011011001000111000) && ({row_reg, col_reg}<18'b011011001000111010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011011001000111010) && ({row_reg, col_reg}<18'b011011001001000000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b011011001001000000)) color_data = 12'b011010101111;
		if(({row_reg, col_reg}>=18'b011011001001000001) && ({row_reg, col_reg}<18'b011011001001011010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011011001001011010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011011001001011011) && ({row_reg, col_reg}<18'b011011001001100111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011011001001100111) && ({row_reg, col_reg}<18'b011011001001101010)) color_data = 12'b011010101111;

		if(({row_reg, col_reg}>=18'b011011001001101010) && ({row_reg, col_reg}<18'b011011010000101110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011011010000101110) && ({row_reg, col_reg}<18'b011011010000110000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011011010000110000) && ({row_reg, col_reg}<18'b011011010000110111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011011010000110111)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011011010000111000) && ({row_reg, col_reg}<18'b011011010000111010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011011010000111010) && ({row_reg, col_reg}<18'b011011010000111100)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011011010000111100) && ({row_reg, col_reg}<18'b011011010001000000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011011010001000000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011011010001000001) && ({row_reg, col_reg}<18'b011011010001001110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011011010001001110) && ({row_reg, col_reg}<18'b011011010001010000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b011011010001010000)) color_data = 12'b011010111110;
		if(({row_reg, col_reg}>=18'b011011010001010001) && ({row_reg, col_reg}<18'b011011010001100100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011011010001100100) && ({row_reg, col_reg}<18'b011011010001110000)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b011011010001110000) && ({row_reg, col_reg}<18'b011011011000101100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011011011000101100) && ({row_reg, col_reg}<18'b011011011000110000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011011011000110000) && ({row_reg, col_reg}<18'b011011011000111001)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011011011000111001) && ({row_reg, col_reg}<18'b011011011000111100)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011011011000111100) && ({row_reg, col_reg}<18'b011011011000111111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011011011000111111) && ({row_reg, col_reg}<18'b011011011001000001)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011011011001000001) && ({row_reg, col_reg}<18'b011011011001000101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011011011001000101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011011011001000110) && ({row_reg, col_reg}<18'b011011011001100110)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011011011001100110) && ({row_reg, col_reg}<18'b011011011001110000)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b011011011001110000) && ({row_reg, col_reg}<18'b011011100001000000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011011100001000000) && ({row_reg, col_reg}<18'b011011100001000110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011011100001000110) && ({row_reg, col_reg}<18'b011011100001100101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011011100001100101) && ({row_reg, col_reg}<18'b011011100001110010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011011100001110010) && ({row_reg, col_reg}<18'b011011100001111111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011011100001111111)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b011011100010000000) && ({row_reg, col_reg}<18'b011011101000110000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011011101000110000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011011101000110001) && ({row_reg, col_reg}<18'b011011101000110011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011011101000110011) && ({row_reg, col_reg}<18'b011011101000110101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011011101000110101) && ({row_reg, col_reg}<18'b011011101000110111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011011101000110111) && ({row_reg, col_reg}<18'b011011101000111001)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011011101000111001) && ({row_reg, col_reg}<18'b011011101000111100)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011011101000111100) && ({row_reg, col_reg}<18'b011011101000111110)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011011101000111110) && ({row_reg, col_reg}<18'b011011101001000000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011011101001000000) && ({row_reg, col_reg}<18'b011011101001000111)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011011101001000111) && ({row_reg, col_reg}<18'b011011101001010010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011011101001010010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011011101001010011) && ({row_reg, col_reg}<18'b011011101001011010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011011101001011010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011011101001011011) && ({row_reg, col_reg}<18'b011011101001100101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011011101001100101) && ({row_reg, col_reg}<18'b011011101001101101)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b011011101001101101) && ({row_reg, col_reg}<18'b011011110000111011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011011110000111011)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011011110000111100) && ({row_reg, col_reg}<18'b011011110001000000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011011110001000000) && ({row_reg, col_reg}<18'b011011110001001000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011011110001001000) && ({row_reg, col_reg}<18'b011011110001010000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011011110001010000) && ({row_reg, col_reg}<18'b011011110001010010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011011110001010010) && ({row_reg, col_reg}<18'b011011110001100101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011011110001100101) && ({row_reg, col_reg}<18'b011011110001101011)) color_data = 12'b011110101110;

		if(({row_reg, col_reg}>=18'b011011110001101011) && ({row_reg, col_reg}<18'b011011111000110000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011011111000110000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011011111000110001) && ({row_reg, col_reg}<18'b011011111000110011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011011111000110011) && ({row_reg, col_reg}<18'b011011111000110101)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011011111000110101) && ({row_reg, col_reg}<18'b011011111000110111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011011111000110111)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011011111000111000) && ({row_reg, col_reg}<18'b011011111000111010)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011011111000111010)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011011111000111011) && ({row_reg, col_reg}<18'b011011111000111111)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011011111000111111) && ({row_reg, col_reg}<18'b011011111001001000)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011011111001001000) && ({row_reg, col_reg}<18'b011011111001010000)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011011111001010000) && ({row_reg, col_reg}<18'b011011111001010011)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}==18'b011011111001010011)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}==18'b011011111001010100)) color_data = 12'b011110101110;
		if(({row_reg, col_reg}>=18'b011011111001010101) && ({row_reg, col_reg}<18'b011011111001100101)) color_data = 12'b011010101110;
		if(({row_reg, col_reg}>=18'b011011111001100101) && ({row_reg, col_reg}<18'b011011111001101010)) color_data = 12'b011110101110;




















































		if(({row_reg, col_reg}>=18'b011011111001101010) && ({row_reg, col_reg}<=18'b100010010100010010)) color_data = 12'b011010101110;
	end
endmodule